// This is the unpowered netlist.
module vga_m (clk_i,
    enable_i,
    fb_i,
    hsync_o,
    nrst_i,
    vsync_o,
    base_h_active_i,
    base_h_bporch_i,
    base_h_fporch_i,
    base_h_sync_i,
    base_v_active_i,
    base_v_bporch_i,
    base_v_fporch_i,
    base_v_sync_i,
    mport_i,
    mport_o,
    pixel_o,
    prescaler_i,
    resolution_i);
 input clk_i;
 input enable_i;
 input fb_i;
 output hsync_o;
 input nrst_i;
 output vsync_o;
 input [9:0] base_h_active_i;
 input [6:0] base_h_bporch_i;
 input [4:0] base_h_fporch_i;
 input [6:0] base_h_sync_i;
 input [8:0] base_v_active_i;
 input [3:0] base_v_bporch_i;
 input [2:0] base_v_fporch_i;
 input [2:0] base_v_sync_i;
 input [33:0] mport_i;
 output [68:0] mport_o;
 output [7:0] pixel_o;
 input [3:0] prescaler_i;
 input [3:0] resolution_i;

 wire net354;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net355;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net356;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net357;
 wire net358;
 wire net359;
 wire net388;
 wire net389;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire \base_h_active[0] ;
 wire \base_h_active[1] ;
 wire \base_h_active[2] ;
 wire \base_h_active[3] ;
 wire \base_h_active[4] ;
 wire \base_h_active[5] ;
 wire \base_h_active[6] ;
 wire \base_h_active[7] ;
 wire \base_h_active[8] ;
 wire \base_h_active[9] ;
 wire \base_h_bporch[0] ;
 wire \base_h_bporch[1] ;
 wire \base_h_bporch[2] ;
 wire \base_h_bporch[3] ;
 wire \base_h_bporch[4] ;
 wire \base_h_bporch[5] ;
 wire \base_h_bporch[6] ;
 wire \base_h_counter[0] ;
 wire \base_h_counter[1] ;
 wire \base_h_counter[2] ;
 wire \base_h_counter[3] ;
 wire \base_h_counter[4] ;
 wire \base_h_counter[5] ;
 wire \base_h_counter[6] ;
 wire \base_h_counter[7] ;
 wire \base_h_counter[8] ;
 wire \base_h_counter[9] ;
 wire \base_h_fporch[0] ;
 wire \base_h_fporch[1] ;
 wire \base_h_fporch[2] ;
 wire \base_h_fporch[3] ;
 wire \base_h_fporch[4] ;
 wire \base_h_sync[0] ;
 wire \base_h_sync[1] ;
 wire \base_h_sync[2] ;
 wire \base_h_sync[3] ;
 wire \base_h_sync[4] ;
 wire \base_h_sync[5] ;
 wire \base_h_sync[6] ;
 wire \base_v_active[0] ;
 wire \base_v_active[1] ;
 wire \base_v_active[2] ;
 wire \base_v_active[3] ;
 wire \base_v_active[4] ;
 wire \base_v_active[5] ;
 wire \base_v_active[6] ;
 wire \base_v_active[7] ;
 wire \base_v_active[8] ;
 wire \base_v_bporch[0] ;
 wire \base_v_bporch[1] ;
 wire \base_v_bporch[2] ;
 wire \base_v_bporch[3] ;
 wire \base_v_counter[0] ;
 wire \base_v_counter[1] ;
 wire \base_v_counter[2] ;
 wire \base_v_counter[3] ;
 wire \base_v_counter[4] ;
 wire \base_v_counter[5] ;
 wire \base_v_counter[6] ;
 wire \base_v_counter[7] ;
 wire \base_v_counter[8] ;
 wire \base_v_counter[9] ;
 wire \base_v_fporch[0] ;
 wire \base_v_fporch[1] ;
 wire \base_v_fporch[2] ;
 wire \base_v_sync[0] ;
 wire \base_v_sync[1] ;
 wire \base_v_sync[2] ;
 wire clknet_0_clk_i;
 wire clknet_2_0_0_clk_i;
 wire clknet_2_1_0_clk_i;
 wire clknet_2_2_0_clk_i;
 wire clknet_2_3_0_clk_i;
 wire clknet_5_0__leaf_clk_i;
 wire clknet_5_10__leaf_clk_i;
 wire clknet_5_11__leaf_clk_i;
 wire clknet_5_12__leaf_clk_i;
 wire clknet_5_13__leaf_clk_i;
 wire clknet_5_14__leaf_clk_i;
 wire clknet_5_15__leaf_clk_i;
 wire clknet_5_16__leaf_clk_i;
 wire clknet_5_17__leaf_clk_i;
 wire clknet_5_18__leaf_clk_i;
 wire clknet_5_19__leaf_clk_i;
 wire clknet_5_1__leaf_clk_i;
 wire clknet_5_20__leaf_clk_i;
 wire clknet_5_21__leaf_clk_i;
 wire clknet_5_22__leaf_clk_i;
 wire clknet_5_23__leaf_clk_i;
 wire clknet_5_24__leaf_clk_i;
 wire clknet_5_25__leaf_clk_i;
 wire clknet_5_26__leaf_clk_i;
 wire clknet_5_27__leaf_clk_i;
 wire clknet_5_28__leaf_clk_i;
 wire clknet_5_29__leaf_clk_i;
 wire clknet_5_2__leaf_clk_i;
 wire clknet_5_30__leaf_clk_i;
 wire clknet_5_31__leaf_clk_i;
 wire clknet_5_3__leaf_clk_i;
 wire clknet_5_4__leaf_clk_i;
 wire clknet_5_5__leaf_clk_i;
 wire clknet_5_6__leaf_clk_i;
 wire clknet_5_7__leaf_clk_i;
 wire clknet_5_8__leaf_clk_i;
 wire clknet_5_9__leaf_clk_i;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_leaf_105_clk_i;
 wire clknet_leaf_106_clk_i;
 wire clknet_leaf_107_clk_i;
 wire clknet_leaf_108_clk_i;
 wire clknet_leaf_109_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_110_clk_i;
 wire clknet_leaf_111_clk_i;
 wire clknet_leaf_112_clk_i;
 wire clknet_leaf_113_clk_i;
 wire clknet_leaf_114_clk_i;
 wire clknet_leaf_115_clk_i;
 wire clknet_leaf_116_clk_i;
 wire clknet_leaf_117_clk_i;
 wire clknet_leaf_118_clk_i;
 wire clknet_leaf_119_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_120_clk_i;
 wire clknet_leaf_121_clk_i;
 wire clknet_leaf_122_clk_i;
 wire clknet_leaf_123_clk_i;
 wire clknet_leaf_124_clk_i;
 wire clknet_leaf_125_clk_i;
 wire clknet_leaf_126_clk_i;
 wire clknet_leaf_127_clk_i;
 wire clknet_leaf_128_clk_i;
 wire clknet_leaf_129_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_130_clk_i;
 wire clknet_leaf_131_clk_i;
 wire clknet_leaf_132_clk_i;
 wire clknet_leaf_133_clk_i;
 wire clknet_leaf_134_clk_i;
 wire clknet_leaf_135_clk_i;
 wire clknet_leaf_136_clk_i;
 wire clknet_leaf_137_clk_i;
 wire clknet_leaf_138_clk_i;
 wire clknet_leaf_139_clk_i;
 wire clknet_leaf_140_clk_i;
 wire clknet_leaf_141_clk_i;
 wire clknet_leaf_142_clk_i;
 wire clknet_leaf_143_clk_i;
 wire clknet_leaf_144_clk_i;
 wire clknet_leaf_145_clk_i;
 wire clknet_leaf_146_clk_i;
 wire clknet_leaf_147_clk_i;
 wire clknet_leaf_148_clk_i;
 wire clknet_leaf_149_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_150_clk_i;
 wire clknet_leaf_151_clk_i;
 wire clknet_leaf_152_clk_i;
 wire clknet_leaf_153_clk_i;
 wire clknet_leaf_154_clk_i;
 wire clknet_leaf_155_clk_i;
 wire clknet_leaf_156_clk_i;
 wire clknet_leaf_157_clk_i;
 wire clknet_leaf_158_clk_i;
 wire clknet_leaf_159_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_160_clk_i;
 wire clknet_leaf_161_clk_i;
 wire clknet_leaf_162_clk_i;
 wire clknet_leaf_163_clk_i;
 wire clknet_leaf_164_clk_i;
 wire clknet_leaf_165_clk_i;
 wire clknet_leaf_166_clk_i;
 wire clknet_leaf_167_clk_i;
 wire clknet_leaf_168_clk_i;
 wire clknet_leaf_169_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_170_clk_i;
 wire clknet_leaf_171_clk_i;
 wire clknet_leaf_172_clk_i;
 wire clknet_leaf_173_clk_i;
 wire clknet_leaf_174_clk_i;
 wire clknet_leaf_175_clk_i;
 wire clknet_leaf_176_clk_i;
 wire clknet_leaf_177_clk_i;
 wire clknet_leaf_178_clk_i;
 wire clknet_leaf_179_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_180_clk_i;
 wire clknet_leaf_181_clk_i;
 wire clknet_leaf_182_clk_i;
 wire clknet_leaf_183_clk_i;
 wire clknet_leaf_184_clk_i;
 wire clknet_leaf_185_clk_i;
 wire clknet_leaf_186_clk_i;
 wire clknet_leaf_187_clk_i;
 wire clknet_leaf_188_clk_i;
 wire clknet_leaf_189_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_190_clk_i;
 wire clknet_leaf_191_clk_i;
 wire clknet_leaf_192_clk_i;
 wire clknet_leaf_193_clk_i;
 wire clknet_leaf_194_clk_i;
 wire clknet_leaf_195_clk_i;
 wire clknet_leaf_196_clk_i;
 wire clknet_leaf_197_clk_i;
 wire clknet_leaf_198_clk_i;
 wire clknet_leaf_199_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_200_clk_i;
 wire clknet_leaf_201_clk_i;
 wire clknet_leaf_202_clk_i;
 wire clknet_leaf_203_clk_i;
 wire clknet_leaf_204_clk_i;
 wire clknet_leaf_205_clk_i;
 wire clknet_leaf_206_clk_i;
 wire clknet_leaf_207_clk_i;
 wire clknet_leaf_208_clk_i;
 wire clknet_leaf_209_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_210_clk_i;
 wire clknet_leaf_211_clk_i;
 wire clknet_leaf_212_clk_i;
 wire clknet_leaf_213_clk_i;
 wire clknet_leaf_214_clk_i;
 wire clknet_leaf_215_clk_i;
 wire clknet_leaf_216_clk_i;
 wire clknet_leaf_217_clk_i;
 wire clknet_leaf_218_clk_i;
 wire clknet_leaf_219_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_220_clk_i;
 wire clknet_leaf_221_clk_i;
 wire clknet_leaf_222_clk_i;
 wire clknet_leaf_223_clk_i;
 wire clknet_leaf_224_clk_i;
 wire clknet_leaf_225_clk_i;
 wire clknet_leaf_226_clk_i;
 wire clknet_leaf_227_clk_i;
 wire clknet_leaf_228_clk_i;
 wire clknet_leaf_229_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_230_clk_i;
 wire clknet_leaf_231_clk_i;
 wire clknet_leaf_232_clk_i;
 wire clknet_leaf_233_clk_i;
 wire clknet_leaf_234_clk_i;
 wire clknet_leaf_235_clk_i;
 wire clknet_leaf_236_clk_i;
 wire clknet_leaf_237_clk_i;
 wire clknet_leaf_238_clk_i;
 wire clknet_leaf_239_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_240_clk_i;
 wire clknet_leaf_241_clk_i;
 wire clknet_leaf_242_clk_i;
 wire clknet_leaf_243_clk_i;
 wire clknet_leaf_244_clk_i;
 wire clknet_leaf_245_clk_i;
 wire clknet_leaf_246_clk_i;
 wire clknet_leaf_247_clk_i;
 wire clknet_leaf_248_clk_i;
 wire clknet_leaf_249_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_250_clk_i;
 wire clknet_leaf_251_clk_i;
 wire clknet_leaf_252_clk_i;
 wire clknet_leaf_253_clk_i;
 wire clknet_leaf_254_clk_i;
 wire clknet_leaf_255_clk_i;
 wire clknet_leaf_256_clk_i;
 wire clknet_leaf_257_clk_i;
 wire clknet_leaf_258_clk_i;
 wire clknet_leaf_259_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_260_clk_i;
 wire clknet_leaf_261_clk_i;
 wire clknet_leaf_262_clk_i;
 wire clknet_leaf_263_clk_i;
 wire clknet_leaf_264_clk_i;
 wire clknet_leaf_265_clk_i;
 wire clknet_leaf_266_clk_i;
 wire clknet_leaf_267_clk_i;
 wire clknet_leaf_268_clk_i;
 wire clknet_leaf_269_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_270_clk_i;
 wire clknet_leaf_271_clk_i;
 wire clknet_leaf_272_clk_i;
 wire clknet_leaf_273_clk_i;
 wire clknet_leaf_274_clk_i;
 wire clknet_leaf_275_clk_i;
 wire clknet_leaf_276_clk_i;
 wire clknet_leaf_277_clk_i;
 wire clknet_leaf_278_clk_i;
 wire clknet_leaf_279_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_280_clk_i;
 wire clknet_leaf_281_clk_i;
 wire clknet_leaf_282_clk_i;
 wire clknet_leaf_283_clk_i;
 wire clknet_leaf_284_clk_i;
 wire clknet_leaf_285_clk_i;
 wire clknet_leaf_286_clk_i;
 wire clknet_leaf_287_clk_i;
 wire clknet_leaf_288_clk_i;
 wire clknet_leaf_289_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_290_clk_i;
 wire clknet_leaf_291_clk_i;
 wire clknet_leaf_292_clk_i;
 wire clknet_leaf_293_clk_i;
 wire clknet_leaf_294_clk_i;
 wire clknet_leaf_295_clk_i;
 wire clknet_leaf_296_clk_i;
 wire clknet_leaf_297_clk_i;
 wire clknet_leaf_298_clk_i;
 wire clknet_leaf_299_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_300_clk_i;
 wire clknet_leaf_301_clk_i;
 wire clknet_leaf_302_clk_i;
 wire clknet_leaf_303_clk_i;
 wire clknet_leaf_304_clk_i;
 wire clknet_leaf_305_clk_i;
 wire clknet_leaf_306_clk_i;
 wire clknet_leaf_307_clk_i;
 wire clknet_leaf_308_clk_i;
 wire clknet_leaf_309_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_310_clk_i;
 wire clknet_leaf_311_clk_i;
 wire clknet_leaf_312_clk_i;
 wire clknet_leaf_313_clk_i;
 wire clknet_leaf_314_clk_i;
 wire clknet_leaf_315_clk_i;
 wire clknet_leaf_316_clk_i;
 wire clknet_leaf_317_clk_i;
 wire clknet_leaf_318_clk_i;
 wire clknet_leaf_319_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_320_clk_i;
 wire clknet_leaf_321_clk_i;
 wire clknet_leaf_322_clk_i;
 wire clknet_leaf_323_clk_i;
 wire clknet_leaf_324_clk_i;
 wire clknet_leaf_325_clk_i;
 wire clknet_leaf_326_clk_i;
 wire clknet_leaf_327_clk_i;
 wire clknet_leaf_328_clk_i;
 wire clknet_leaf_329_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_330_clk_i;
 wire clknet_leaf_331_clk_i;
 wire clknet_leaf_332_clk_i;
 wire clknet_leaf_333_clk_i;
 wire clknet_leaf_334_clk_i;
 wire clknet_leaf_335_clk_i;
 wire clknet_leaf_336_clk_i;
 wire clknet_leaf_337_clk_i;
 wire clknet_leaf_338_clk_i;
 wire clknet_leaf_339_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_340_clk_i;
 wire clknet_leaf_341_clk_i;
 wire clknet_leaf_342_clk_i;
 wire clknet_leaf_343_clk_i;
 wire clknet_leaf_344_clk_i;
 wire clknet_leaf_345_clk_i;
 wire clknet_leaf_346_clk_i;
 wire clknet_leaf_347_clk_i;
 wire clknet_leaf_348_clk_i;
 wire clknet_leaf_349_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_350_clk_i;
 wire clknet_leaf_351_clk_i;
 wire clknet_leaf_352_clk_i;
 wire clknet_leaf_353_clk_i;
 wire clknet_leaf_354_clk_i;
 wire clknet_leaf_355_clk_i;
 wire clknet_leaf_356_clk_i;
 wire clknet_leaf_357_clk_i;
 wire clknet_leaf_358_clk_i;
 wire clknet_leaf_359_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_360_clk_i;
 wire clknet_leaf_361_clk_i;
 wire clknet_leaf_362_clk_i;
 wire clknet_leaf_363_clk_i;
 wire clknet_leaf_364_clk_i;
 wire clknet_leaf_365_clk_i;
 wire clknet_leaf_366_clk_i;
 wire clknet_leaf_367_clk_i;
 wire clknet_leaf_368_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_370_clk_i;
 wire clknet_leaf_371_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_46_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_50_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_54_clk_i;
 wire clknet_leaf_55_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_58_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_62_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_65_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_68_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_72_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_76_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_80_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_82_clk_i;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_84_clk_i;
 wire clknet_leaf_85_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_90_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_9_clk_i;
 wire \fb_read_state[0] ;
 wire \fb_read_state[1] ;
 wire \fb_read_state[2] ;
 wire \line_cache[0][0] ;
 wire \line_cache[0][1] ;
 wire \line_cache[0][2] ;
 wire \line_cache[0][3] ;
 wire \line_cache[0][4] ;
 wire \line_cache[0][5] ;
 wire \line_cache[0][6] ;
 wire \line_cache[0][7] ;
 wire \line_cache[100][0] ;
 wire \line_cache[100][1] ;
 wire \line_cache[100][2] ;
 wire \line_cache[100][3] ;
 wire \line_cache[100][4] ;
 wire \line_cache[100][5] ;
 wire \line_cache[100][6] ;
 wire \line_cache[100][7] ;
 wire \line_cache[101][0] ;
 wire \line_cache[101][1] ;
 wire \line_cache[101][2] ;
 wire \line_cache[101][3] ;
 wire \line_cache[101][4] ;
 wire \line_cache[101][5] ;
 wire \line_cache[101][6] ;
 wire \line_cache[101][7] ;
 wire \line_cache[102][0] ;
 wire \line_cache[102][1] ;
 wire \line_cache[102][2] ;
 wire \line_cache[102][3] ;
 wire \line_cache[102][4] ;
 wire \line_cache[102][5] ;
 wire \line_cache[102][6] ;
 wire \line_cache[102][7] ;
 wire \line_cache[103][0] ;
 wire \line_cache[103][1] ;
 wire \line_cache[103][2] ;
 wire \line_cache[103][3] ;
 wire \line_cache[103][4] ;
 wire \line_cache[103][5] ;
 wire \line_cache[103][6] ;
 wire \line_cache[103][7] ;
 wire \line_cache[104][0] ;
 wire \line_cache[104][1] ;
 wire \line_cache[104][2] ;
 wire \line_cache[104][3] ;
 wire \line_cache[104][4] ;
 wire \line_cache[104][5] ;
 wire \line_cache[104][6] ;
 wire \line_cache[104][7] ;
 wire \line_cache[105][0] ;
 wire \line_cache[105][1] ;
 wire \line_cache[105][2] ;
 wire \line_cache[105][3] ;
 wire \line_cache[105][4] ;
 wire \line_cache[105][5] ;
 wire \line_cache[105][6] ;
 wire \line_cache[105][7] ;
 wire \line_cache[106][0] ;
 wire \line_cache[106][1] ;
 wire \line_cache[106][2] ;
 wire \line_cache[106][3] ;
 wire \line_cache[106][4] ;
 wire \line_cache[106][5] ;
 wire \line_cache[106][6] ;
 wire \line_cache[106][7] ;
 wire \line_cache[107][0] ;
 wire \line_cache[107][1] ;
 wire \line_cache[107][2] ;
 wire \line_cache[107][3] ;
 wire \line_cache[107][4] ;
 wire \line_cache[107][5] ;
 wire \line_cache[107][6] ;
 wire \line_cache[107][7] ;
 wire \line_cache[108][0] ;
 wire \line_cache[108][1] ;
 wire \line_cache[108][2] ;
 wire \line_cache[108][3] ;
 wire \line_cache[108][4] ;
 wire \line_cache[108][5] ;
 wire \line_cache[108][6] ;
 wire \line_cache[108][7] ;
 wire \line_cache[109][0] ;
 wire \line_cache[109][1] ;
 wire \line_cache[109][2] ;
 wire \line_cache[109][3] ;
 wire \line_cache[109][4] ;
 wire \line_cache[109][5] ;
 wire \line_cache[109][6] ;
 wire \line_cache[109][7] ;
 wire \line_cache[10][0] ;
 wire \line_cache[10][1] ;
 wire \line_cache[10][2] ;
 wire \line_cache[10][3] ;
 wire \line_cache[10][4] ;
 wire \line_cache[10][5] ;
 wire \line_cache[10][6] ;
 wire \line_cache[10][7] ;
 wire \line_cache[110][0] ;
 wire \line_cache[110][1] ;
 wire \line_cache[110][2] ;
 wire \line_cache[110][3] ;
 wire \line_cache[110][4] ;
 wire \line_cache[110][5] ;
 wire \line_cache[110][6] ;
 wire \line_cache[110][7] ;
 wire \line_cache[111][0] ;
 wire \line_cache[111][1] ;
 wire \line_cache[111][2] ;
 wire \line_cache[111][3] ;
 wire \line_cache[111][4] ;
 wire \line_cache[111][5] ;
 wire \line_cache[111][6] ;
 wire \line_cache[111][7] ;
 wire \line_cache[112][0] ;
 wire \line_cache[112][1] ;
 wire \line_cache[112][2] ;
 wire \line_cache[112][3] ;
 wire \line_cache[112][4] ;
 wire \line_cache[112][5] ;
 wire \line_cache[112][6] ;
 wire \line_cache[112][7] ;
 wire \line_cache[113][0] ;
 wire \line_cache[113][1] ;
 wire \line_cache[113][2] ;
 wire \line_cache[113][3] ;
 wire \line_cache[113][4] ;
 wire \line_cache[113][5] ;
 wire \line_cache[113][6] ;
 wire \line_cache[113][7] ;
 wire \line_cache[114][0] ;
 wire \line_cache[114][1] ;
 wire \line_cache[114][2] ;
 wire \line_cache[114][3] ;
 wire \line_cache[114][4] ;
 wire \line_cache[114][5] ;
 wire \line_cache[114][6] ;
 wire \line_cache[114][7] ;
 wire \line_cache[115][0] ;
 wire \line_cache[115][1] ;
 wire \line_cache[115][2] ;
 wire \line_cache[115][3] ;
 wire \line_cache[115][4] ;
 wire \line_cache[115][5] ;
 wire \line_cache[115][6] ;
 wire \line_cache[115][7] ;
 wire \line_cache[116][0] ;
 wire \line_cache[116][1] ;
 wire \line_cache[116][2] ;
 wire \line_cache[116][3] ;
 wire \line_cache[116][4] ;
 wire \line_cache[116][5] ;
 wire \line_cache[116][6] ;
 wire \line_cache[116][7] ;
 wire \line_cache[117][0] ;
 wire \line_cache[117][1] ;
 wire \line_cache[117][2] ;
 wire \line_cache[117][3] ;
 wire \line_cache[117][4] ;
 wire \line_cache[117][5] ;
 wire \line_cache[117][6] ;
 wire \line_cache[117][7] ;
 wire \line_cache[118][0] ;
 wire \line_cache[118][1] ;
 wire \line_cache[118][2] ;
 wire \line_cache[118][3] ;
 wire \line_cache[118][4] ;
 wire \line_cache[118][5] ;
 wire \line_cache[118][6] ;
 wire \line_cache[118][7] ;
 wire \line_cache[119][0] ;
 wire \line_cache[119][1] ;
 wire \line_cache[119][2] ;
 wire \line_cache[119][3] ;
 wire \line_cache[119][4] ;
 wire \line_cache[119][5] ;
 wire \line_cache[119][6] ;
 wire \line_cache[119][7] ;
 wire \line_cache[11][0] ;
 wire \line_cache[11][1] ;
 wire \line_cache[11][2] ;
 wire \line_cache[11][3] ;
 wire \line_cache[11][4] ;
 wire \line_cache[11][5] ;
 wire \line_cache[11][6] ;
 wire \line_cache[11][7] ;
 wire \line_cache[120][0] ;
 wire \line_cache[120][1] ;
 wire \line_cache[120][2] ;
 wire \line_cache[120][3] ;
 wire \line_cache[120][4] ;
 wire \line_cache[120][5] ;
 wire \line_cache[120][6] ;
 wire \line_cache[120][7] ;
 wire \line_cache[121][0] ;
 wire \line_cache[121][1] ;
 wire \line_cache[121][2] ;
 wire \line_cache[121][3] ;
 wire \line_cache[121][4] ;
 wire \line_cache[121][5] ;
 wire \line_cache[121][6] ;
 wire \line_cache[121][7] ;
 wire \line_cache[122][0] ;
 wire \line_cache[122][1] ;
 wire \line_cache[122][2] ;
 wire \line_cache[122][3] ;
 wire \line_cache[122][4] ;
 wire \line_cache[122][5] ;
 wire \line_cache[122][6] ;
 wire \line_cache[122][7] ;
 wire \line_cache[123][0] ;
 wire \line_cache[123][1] ;
 wire \line_cache[123][2] ;
 wire \line_cache[123][3] ;
 wire \line_cache[123][4] ;
 wire \line_cache[123][5] ;
 wire \line_cache[123][6] ;
 wire \line_cache[123][7] ;
 wire \line_cache[124][0] ;
 wire \line_cache[124][1] ;
 wire \line_cache[124][2] ;
 wire \line_cache[124][3] ;
 wire \line_cache[124][4] ;
 wire \line_cache[124][5] ;
 wire \line_cache[124][6] ;
 wire \line_cache[124][7] ;
 wire \line_cache[125][0] ;
 wire \line_cache[125][1] ;
 wire \line_cache[125][2] ;
 wire \line_cache[125][3] ;
 wire \line_cache[125][4] ;
 wire \line_cache[125][5] ;
 wire \line_cache[125][6] ;
 wire \line_cache[125][7] ;
 wire \line_cache[126][0] ;
 wire \line_cache[126][1] ;
 wire \line_cache[126][2] ;
 wire \line_cache[126][3] ;
 wire \line_cache[126][4] ;
 wire \line_cache[126][5] ;
 wire \line_cache[126][6] ;
 wire \line_cache[126][7] ;
 wire \line_cache[127][0] ;
 wire \line_cache[127][1] ;
 wire \line_cache[127][2] ;
 wire \line_cache[127][3] ;
 wire \line_cache[127][4] ;
 wire \line_cache[127][5] ;
 wire \line_cache[127][6] ;
 wire \line_cache[127][7] ;
 wire \line_cache[128][0] ;
 wire \line_cache[128][1] ;
 wire \line_cache[128][2] ;
 wire \line_cache[128][3] ;
 wire \line_cache[128][4] ;
 wire \line_cache[128][5] ;
 wire \line_cache[128][6] ;
 wire \line_cache[128][7] ;
 wire \line_cache[129][0] ;
 wire \line_cache[129][1] ;
 wire \line_cache[129][2] ;
 wire \line_cache[129][3] ;
 wire \line_cache[129][4] ;
 wire \line_cache[129][5] ;
 wire \line_cache[129][6] ;
 wire \line_cache[129][7] ;
 wire \line_cache[12][0] ;
 wire \line_cache[12][1] ;
 wire \line_cache[12][2] ;
 wire \line_cache[12][3] ;
 wire \line_cache[12][4] ;
 wire \line_cache[12][5] ;
 wire \line_cache[12][6] ;
 wire \line_cache[12][7] ;
 wire \line_cache[130][0] ;
 wire \line_cache[130][1] ;
 wire \line_cache[130][2] ;
 wire \line_cache[130][3] ;
 wire \line_cache[130][4] ;
 wire \line_cache[130][5] ;
 wire \line_cache[130][6] ;
 wire \line_cache[130][7] ;
 wire \line_cache[131][0] ;
 wire \line_cache[131][1] ;
 wire \line_cache[131][2] ;
 wire \line_cache[131][3] ;
 wire \line_cache[131][4] ;
 wire \line_cache[131][5] ;
 wire \line_cache[131][6] ;
 wire \line_cache[131][7] ;
 wire \line_cache[132][0] ;
 wire \line_cache[132][1] ;
 wire \line_cache[132][2] ;
 wire \line_cache[132][3] ;
 wire \line_cache[132][4] ;
 wire \line_cache[132][5] ;
 wire \line_cache[132][6] ;
 wire \line_cache[132][7] ;
 wire \line_cache[133][0] ;
 wire \line_cache[133][1] ;
 wire \line_cache[133][2] ;
 wire \line_cache[133][3] ;
 wire \line_cache[133][4] ;
 wire \line_cache[133][5] ;
 wire \line_cache[133][6] ;
 wire \line_cache[133][7] ;
 wire \line_cache[134][0] ;
 wire \line_cache[134][1] ;
 wire \line_cache[134][2] ;
 wire \line_cache[134][3] ;
 wire \line_cache[134][4] ;
 wire \line_cache[134][5] ;
 wire \line_cache[134][6] ;
 wire \line_cache[134][7] ;
 wire \line_cache[135][0] ;
 wire \line_cache[135][1] ;
 wire \line_cache[135][2] ;
 wire \line_cache[135][3] ;
 wire \line_cache[135][4] ;
 wire \line_cache[135][5] ;
 wire \line_cache[135][6] ;
 wire \line_cache[135][7] ;
 wire \line_cache[136][0] ;
 wire \line_cache[136][1] ;
 wire \line_cache[136][2] ;
 wire \line_cache[136][3] ;
 wire \line_cache[136][4] ;
 wire \line_cache[136][5] ;
 wire \line_cache[136][6] ;
 wire \line_cache[136][7] ;
 wire \line_cache[137][0] ;
 wire \line_cache[137][1] ;
 wire \line_cache[137][2] ;
 wire \line_cache[137][3] ;
 wire \line_cache[137][4] ;
 wire \line_cache[137][5] ;
 wire \line_cache[137][6] ;
 wire \line_cache[137][7] ;
 wire \line_cache[138][0] ;
 wire \line_cache[138][1] ;
 wire \line_cache[138][2] ;
 wire \line_cache[138][3] ;
 wire \line_cache[138][4] ;
 wire \line_cache[138][5] ;
 wire \line_cache[138][6] ;
 wire \line_cache[138][7] ;
 wire \line_cache[139][0] ;
 wire \line_cache[139][1] ;
 wire \line_cache[139][2] ;
 wire \line_cache[139][3] ;
 wire \line_cache[139][4] ;
 wire \line_cache[139][5] ;
 wire \line_cache[139][6] ;
 wire \line_cache[139][7] ;
 wire \line_cache[13][0] ;
 wire \line_cache[13][1] ;
 wire \line_cache[13][2] ;
 wire \line_cache[13][3] ;
 wire \line_cache[13][4] ;
 wire \line_cache[13][5] ;
 wire \line_cache[13][6] ;
 wire \line_cache[13][7] ;
 wire \line_cache[140][0] ;
 wire \line_cache[140][1] ;
 wire \line_cache[140][2] ;
 wire \line_cache[140][3] ;
 wire \line_cache[140][4] ;
 wire \line_cache[140][5] ;
 wire \line_cache[140][6] ;
 wire \line_cache[140][7] ;
 wire \line_cache[141][0] ;
 wire \line_cache[141][1] ;
 wire \line_cache[141][2] ;
 wire \line_cache[141][3] ;
 wire \line_cache[141][4] ;
 wire \line_cache[141][5] ;
 wire \line_cache[141][6] ;
 wire \line_cache[141][7] ;
 wire \line_cache[142][0] ;
 wire \line_cache[142][1] ;
 wire \line_cache[142][2] ;
 wire \line_cache[142][3] ;
 wire \line_cache[142][4] ;
 wire \line_cache[142][5] ;
 wire \line_cache[142][6] ;
 wire \line_cache[142][7] ;
 wire \line_cache[143][0] ;
 wire \line_cache[143][1] ;
 wire \line_cache[143][2] ;
 wire \line_cache[143][3] ;
 wire \line_cache[143][4] ;
 wire \line_cache[143][5] ;
 wire \line_cache[143][6] ;
 wire \line_cache[143][7] ;
 wire \line_cache[144][0] ;
 wire \line_cache[144][1] ;
 wire \line_cache[144][2] ;
 wire \line_cache[144][3] ;
 wire \line_cache[144][4] ;
 wire \line_cache[144][5] ;
 wire \line_cache[144][6] ;
 wire \line_cache[144][7] ;
 wire \line_cache[145][0] ;
 wire \line_cache[145][1] ;
 wire \line_cache[145][2] ;
 wire \line_cache[145][3] ;
 wire \line_cache[145][4] ;
 wire \line_cache[145][5] ;
 wire \line_cache[145][6] ;
 wire \line_cache[145][7] ;
 wire \line_cache[146][0] ;
 wire \line_cache[146][1] ;
 wire \line_cache[146][2] ;
 wire \line_cache[146][3] ;
 wire \line_cache[146][4] ;
 wire \line_cache[146][5] ;
 wire \line_cache[146][6] ;
 wire \line_cache[146][7] ;
 wire \line_cache[147][0] ;
 wire \line_cache[147][1] ;
 wire \line_cache[147][2] ;
 wire \line_cache[147][3] ;
 wire \line_cache[147][4] ;
 wire \line_cache[147][5] ;
 wire \line_cache[147][6] ;
 wire \line_cache[147][7] ;
 wire \line_cache[148][0] ;
 wire \line_cache[148][1] ;
 wire \line_cache[148][2] ;
 wire \line_cache[148][3] ;
 wire \line_cache[148][4] ;
 wire \line_cache[148][5] ;
 wire \line_cache[148][6] ;
 wire \line_cache[148][7] ;
 wire \line_cache[149][0] ;
 wire \line_cache[149][1] ;
 wire \line_cache[149][2] ;
 wire \line_cache[149][3] ;
 wire \line_cache[149][4] ;
 wire \line_cache[149][5] ;
 wire \line_cache[149][6] ;
 wire \line_cache[149][7] ;
 wire \line_cache[14][0] ;
 wire \line_cache[14][1] ;
 wire \line_cache[14][2] ;
 wire \line_cache[14][3] ;
 wire \line_cache[14][4] ;
 wire \line_cache[14][5] ;
 wire \line_cache[14][6] ;
 wire \line_cache[14][7] ;
 wire \line_cache[150][0] ;
 wire \line_cache[150][1] ;
 wire \line_cache[150][2] ;
 wire \line_cache[150][3] ;
 wire \line_cache[150][4] ;
 wire \line_cache[150][5] ;
 wire \line_cache[150][6] ;
 wire \line_cache[150][7] ;
 wire \line_cache[151][0] ;
 wire \line_cache[151][1] ;
 wire \line_cache[151][2] ;
 wire \line_cache[151][3] ;
 wire \line_cache[151][4] ;
 wire \line_cache[151][5] ;
 wire \line_cache[151][6] ;
 wire \line_cache[151][7] ;
 wire \line_cache[152][0] ;
 wire \line_cache[152][1] ;
 wire \line_cache[152][2] ;
 wire \line_cache[152][3] ;
 wire \line_cache[152][4] ;
 wire \line_cache[152][5] ;
 wire \line_cache[152][6] ;
 wire \line_cache[152][7] ;
 wire \line_cache[153][0] ;
 wire \line_cache[153][1] ;
 wire \line_cache[153][2] ;
 wire \line_cache[153][3] ;
 wire \line_cache[153][4] ;
 wire \line_cache[153][5] ;
 wire \line_cache[153][6] ;
 wire \line_cache[153][7] ;
 wire \line_cache[154][0] ;
 wire \line_cache[154][1] ;
 wire \line_cache[154][2] ;
 wire \line_cache[154][3] ;
 wire \line_cache[154][4] ;
 wire \line_cache[154][5] ;
 wire \line_cache[154][6] ;
 wire \line_cache[154][7] ;
 wire \line_cache[155][0] ;
 wire \line_cache[155][1] ;
 wire \line_cache[155][2] ;
 wire \line_cache[155][3] ;
 wire \line_cache[155][4] ;
 wire \line_cache[155][5] ;
 wire \line_cache[155][6] ;
 wire \line_cache[155][7] ;
 wire \line_cache[156][0] ;
 wire \line_cache[156][1] ;
 wire \line_cache[156][2] ;
 wire \line_cache[156][3] ;
 wire \line_cache[156][4] ;
 wire \line_cache[156][5] ;
 wire \line_cache[156][6] ;
 wire \line_cache[156][7] ;
 wire \line_cache[157][0] ;
 wire \line_cache[157][1] ;
 wire \line_cache[157][2] ;
 wire \line_cache[157][3] ;
 wire \line_cache[157][4] ;
 wire \line_cache[157][5] ;
 wire \line_cache[157][6] ;
 wire \line_cache[157][7] ;
 wire \line_cache[158][0] ;
 wire \line_cache[158][1] ;
 wire \line_cache[158][2] ;
 wire \line_cache[158][3] ;
 wire \line_cache[158][4] ;
 wire \line_cache[158][5] ;
 wire \line_cache[158][6] ;
 wire \line_cache[158][7] ;
 wire \line_cache[159][0] ;
 wire \line_cache[159][1] ;
 wire \line_cache[159][2] ;
 wire \line_cache[159][3] ;
 wire \line_cache[159][4] ;
 wire \line_cache[159][5] ;
 wire \line_cache[159][6] ;
 wire \line_cache[159][7] ;
 wire \line_cache[15][0] ;
 wire \line_cache[15][1] ;
 wire \line_cache[15][2] ;
 wire \line_cache[15][3] ;
 wire \line_cache[15][4] ;
 wire \line_cache[15][5] ;
 wire \line_cache[15][6] ;
 wire \line_cache[15][7] ;
 wire \line_cache[160][0] ;
 wire \line_cache[160][1] ;
 wire \line_cache[160][2] ;
 wire \line_cache[160][3] ;
 wire \line_cache[160][4] ;
 wire \line_cache[160][5] ;
 wire \line_cache[160][6] ;
 wire \line_cache[160][7] ;
 wire \line_cache[161][0] ;
 wire \line_cache[161][1] ;
 wire \line_cache[161][2] ;
 wire \line_cache[161][3] ;
 wire \line_cache[161][4] ;
 wire \line_cache[161][5] ;
 wire \line_cache[161][6] ;
 wire \line_cache[161][7] ;
 wire \line_cache[162][0] ;
 wire \line_cache[162][1] ;
 wire \line_cache[162][2] ;
 wire \line_cache[162][3] ;
 wire \line_cache[162][4] ;
 wire \line_cache[162][5] ;
 wire \line_cache[162][6] ;
 wire \line_cache[162][7] ;
 wire \line_cache[163][0] ;
 wire \line_cache[163][1] ;
 wire \line_cache[163][2] ;
 wire \line_cache[163][3] ;
 wire \line_cache[163][4] ;
 wire \line_cache[163][5] ;
 wire \line_cache[163][6] ;
 wire \line_cache[163][7] ;
 wire \line_cache[164][0] ;
 wire \line_cache[164][1] ;
 wire \line_cache[164][2] ;
 wire \line_cache[164][3] ;
 wire \line_cache[164][4] ;
 wire \line_cache[164][5] ;
 wire \line_cache[164][6] ;
 wire \line_cache[164][7] ;
 wire \line_cache[165][0] ;
 wire \line_cache[165][1] ;
 wire \line_cache[165][2] ;
 wire \line_cache[165][3] ;
 wire \line_cache[165][4] ;
 wire \line_cache[165][5] ;
 wire \line_cache[165][6] ;
 wire \line_cache[165][7] ;
 wire \line_cache[166][0] ;
 wire \line_cache[166][1] ;
 wire \line_cache[166][2] ;
 wire \line_cache[166][3] ;
 wire \line_cache[166][4] ;
 wire \line_cache[166][5] ;
 wire \line_cache[166][6] ;
 wire \line_cache[166][7] ;
 wire \line_cache[167][0] ;
 wire \line_cache[167][1] ;
 wire \line_cache[167][2] ;
 wire \line_cache[167][3] ;
 wire \line_cache[167][4] ;
 wire \line_cache[167][5] ;
 wire \line_cache[167][6] ;
 wire \line_cache[167][7] ;
 wire \line_cache[168][0] ;
 wire \line_cache[168][1] ;
 wire \line_cache[168][2] ;
 wire \line_cache[168][3] ;
 wire \line_cache[168][4] ;
 wire \line_cache[168][5] ;
 wire \line_cache[168][6] ;
 wire \line_cache[168][7] ;
 wire \line_cache[169][0] ;
 wire \line_cache[169][1] ;
 wire \line_cache[169][2] ;
 wire \line_cache[169][3] ;
 wire \line_cache[169][4] ;
 wire \line_cache[169][5] ;
 wire \line_cache[169][6] ;
 wire \line_cache[169][7] ;
 wire \line_cache[16][0] ;
 wire \line_cache[16][1] ;
 wire \line_cache[16][2] ;
 wire \line_cache[16][3] ;
 wire \line_cache[16][4] ;
 wire \line_cache[16][5] ;
 wire \line_cache[16][6] ;
 wire \line_cache[16][7] ;
 wire \line_cache[170][0] ;
 wire \line_cache[170][1] ;
 wire \line_cache[170][2] ;
 wire \line_cache[170][3] ;
 wire \line_cache[170][4] ;
 wire \line_cache[170][5] ;
 wire \line_cache[170][6] ;
 wire \line_cache[170][7] ;
 wire \line_cache[171][0] ;
 wire \line_cache[171][1] ;
 wire \line_cache[171][2] ;
 wire \line_cache[171][3] ;
 wire \line_cache[171][4] ;
 wire \line_cache[171][5] ;
 wire \line_cache[171][6] ;
 wire \line_cache[171][7] ;
 wire \line_cache[172][0] ;
 wire \line_cache[172][1] ;
 wire \line_cache[172][2] ;
 wire \line_cache[172][3] ;
 wire \line_cache[172][4] ;
 wire \line_cache[172][5] ;
 wire \line_cache[172][6] ;
 wire \line_cache[172][7] ;
 wire \line_cache[173][0] ;
 wire \line_cache[173][1] ;
 wire \line_cache[173][2] ;
 wire \line_cache[173][3] ;
 wire \line_cache[173][4] ;
 wire \line_cache[173][5] ;
 wire \line_cache[173][6] ;
 wire \line_cache[173][7] ;
 wire \line_cache[174][0] ;
 wire \line_cache[174][1] ;
 wire \line_cache[174][2] ;
 wire \line_cache[174][3] ;
 wire \line_cache[174][4] ;
 wire \line_cache[174][5] ;
 wire \line_cache[174][6] ;
 wire \line_cache[174][7] ;
 wire \line_cache[175][0] ;
 wire \line_cache[175][1] ;
 wire \line_cache[175][2] ;
 wire \line_cache[175][3] ;
 wire \line_cache[175][4] ;
 wire \line_cache[175][5] ;
 wire \line_cache[175][6] ;
 wire \line_cache[175][7] ;
 wire \line_cache[176][0] ;
 wire \line_cache[176][1] ;
 wire \line_cache[176][2] ;
 wire \line_cache[176][3] ;
 wire \line_cache[176][4] ;
 wire \line_cache[176][5] ;
 wire \line_cache[176][6] ;
 wire \line_cache[176][7] ;
 wire \line_cache[177][0] ;
 wire \line_cache[177][1] ;
 wire \line_cache[177][2] ;
 wire \line_cache[177][3] ;
 wire \line_cache[177][4] ;
 wire \line_cache[177][5] ;
 wire \line_cache[177][6] ;
 wire \line_cache[177][7] ;
 wire \line_cache[178][0] ;
 wire \line_cache[178][1] ;
 wire \line_cache[178][2] ;
 wire \line_cache[178][3] ;
 wire \line_cache[178][4] ;
 wire \line_cache[178][5] ;
 wire \line_cache[178][6] ;
 wire \line_cache[178][7] ;
 wire \line_cache[179][0] ;
 wire \line_cache[179][1] ;
 wire \line_cache[179][2] ;
 wire \line_cache[179][3] ;
 wire \line_cache[179][4] ;
 wire \line_cache[179][5] ;
 wire \line_cache[179][6] ;
 wire \line_cache[179][7] ;
 wire \line_cache[17][0] ;
 wire \line_cache[17][1] ;
 wire \line_cache[17][2] ;
 wire \line_cache[17][3] ;
 wire \line_cache[17][4] ;
 wire \line_cache[17][5] ;
 wire \line_cache[17][6] ;
 wire \line_cache[17][7] ;
 wire \line_cache[180][0] ;
 wire \line_cache[180][1] ;
 wire \line_cache[180][2] ;
 wire \line_cache[180][3] ;
 wire \line_cache[180][4] ;
 wire \line_cache[180][5] ;
 wire \line_cache[180][6] ;
 wire \line_cache[180][7] ;
 wire \line_cache[181][0] ;
 wire \line_cache[181][1] ;
 wire \line_cache[181][2] ;
 wire \line_cache[181][3] ;
 wire \line_cache[181][4] ;
 wire \line_cache[181][5] ;
 wire \line_cache[181][6] ;
 wire \line_cache[181][7] ;
 wire \line_cache[182][0] ;
 wire \line_cache[182][1] ;
 wire \line_cache[182][2] ;
 wire \line_cache[182][3] ;
 wire \line_cache[182][4] ;
 wire \line_cache[182][5] ;
 wire \line_cache[182][6] ;
 wire \line_cache[182][7] ;
 wire \line_cache[183][0] ;
 wire \line_cache[183][1] ;
 wire \line_cache[183][2] ;
 wire \line_cache[183][3] ;
 wire \line_cache[183][4] ;
 wire \line_cache[183][5] ;
 wire \line_cache[183][6] ;
 wire \line_cache[183][7] ;
 wire \line_cache[184][0] ;
 wire \line_cache[184][1] ;
 wire \line_cache[184][2] ;
 wire \line_cache[184][3] ;
 wire \line_cache[184][4] ;
 wire \line_cache[184][5] ;
 wire \line_cache[184][6] ;
 wire \line_cache[184][7] ;
 wire \line_cache[185][0] ;
 wire \line_cache[185][1] ;
 wire \line_cache[185][2] ;
 wire \line_cache[185][3] ;
 wire \line_cache[185][4] ;
 wire \line_cache[185][5] ;
 wire \line_cache[185][6] ;
 wire \line_cache[185][7] ;
 wire \line_cache[186][0] ;
 wire \line_cache[186][1] ;
 wire \line_cache[186][2] ;
 wire \line_cache[186][3] ;
 wire \line_cache[186][4] ;
 wire \line_cache[186][5] ;
 wire \line_cache[186][6] ;
 wire \line_cache[186][7] ;
 wire \line_cache[187][0] ;
 wire \line_cache[187][1] ;
 wire \line_cache[187][2] ;
 wire \line_cache[187][3] ;
 wire \line_cache[187][4] ;
 wire \line_cache[187][5] ;
 wire \line_cache[187][6] ;
 wire \line_cache[187][7] ;
 wire \line_cache[188][0] ;
 wire \line_cache[188][1] ;
 wire \line_cache[188][2] ;
 wire \line_cache[188][3] ;
 wire \line_cache[188][4] ;
 wire \line_cache[188][5] ;
 wire \line_cache[188][6] ;
 wire \line_cache[188][7] ;
 wire \line_cache[189][0] ;
 wire \line_cache[189][1] ;
 wire \line_cache[189][2] ;
 wire \line_cache[189][3] ;
 wire \line_cache[189][4] ;
 wire \line_cache[189][5] ;
 wire \line_cache[189][6] ;
 wire \line_cache[189][7] ;
 wire \line_cache[18][0] ;
 wire \line_cache[18][1] ;
 wire \line_cache[18][2] ;
 wire \line_cache[18][3] ;
 wire \line_cache[18][4] ;
 wire \line_cache[18][5] ;
 wire \line_cache[18][6] ;
 wire \line_cache[18][7] ;
 wire \line_cache[190][0] ;
 wire \line_cache[190][1] ;
 wire \line_cache[190][2] ;
 wire \line_cache[190][3] ;
 wire \line_cache[190][4] ;
 wire \line_cache[190][5] ;
 wire \line_cache[190][6] ;
 wire \line_cache[190][7] ;
 wire \line_cache[191][0] ;
 wire \line_cache[191][1] ;
 wire \line_cache[191][2] ;
 wire \line_cache[191][3] ;
 wire \line_cache[191][4] ;
 wire \line_cache[191][5] ;
 wire \line_cache[191][6] ;
 wire \line_cache[191][7] ;
 wire \line_cache[192][0] ;
 wire \line_cache[192][1] ;
 wire \line_cache[192][2] ;
 wire \line_cache[192][3] ;
 wire \line_cache[192][4] ;
 wire \line_cache[192][5] ;
 wire \line_cache[192][6] ;
 wire \line_cache[192][7] ;
 wire \line_cache[193][0] ;
 wire \line_cache[193][1] ;
 wire \line_cache[193][2] ;
 wire \line_cache[193][3] ;
 wire \line_cache[193][4] ;
 wire \line_cache[193][5] ;
 wire \line_cache[193][6] ;
 wire \line_cache[193][7] ;
 wire \line_cache[194][0] ;
 wire \line_cache[194][1] ;
 wire \line_cache[194][2] ;
 wire \line_cache[194][3] ;
 wire \line_cache[194][4] ;
 wire \line_cache[194][5] ;
 wire \line_cache[194][6] ;
 wire \line_cache[194][7] ;
 wire \line_cache[195][0] ;
 wire \line_cache[195][1] ;
 wire \line_cache[195][2] ;
 wire \line_cache[195][3] ;
 wire \line_cache[195][4] ;
 wire \line_cache[195][5] ;
 wire \line_cache[195][6] ;
 wire \line_cache[195][7] ;
 wire \line_cache[196][0] ;
 wire \line_cache[196][1] ;
 wire \line_cache[196][2] ;
 wire \line_cache[196][3] ;
 wire \line_cache[196][4] ;
 wire \line_cache[196][5] ;
 wire \line_cache[196][6] ;
 wire \line_cache[196][7] ;
 wire \line_cache[197][0] ;
 wire \line_cache[197][1] ;
 wire \line_cache[197][2] ;
 wire \line_cache[197][3] ;
 wire \line_cache[197][4] ;
 wire \line_cache[197][5] ;
 wire \line_cache[197][6] ;
 wire \line_cache[197][7] ;
 wire \line_cache[198][0] ;
 wire \line_cache[198][1] ;
 wire \line_cache[198][2] ;
 wire \line_cache[198][3] ;
 wire \line_cache[198][4] ;
 wire \line_cache[198][5] ;
 wire \line_cache[198][6] ;
 wire \line_cache[198][7] ;
 wire \line_cache[199][0] ;
 wire \line_cache[199][1] ;
 wire \line_cache[199][2] ;
 wire \line_cache[199][3] ;
 wire \line_cache[199][4] ;
 wire \line_cache[199][5] ;
 wire \line_cache[199][6] ;
 wire \line_cache[199][7] ;
 wire \line_cache[19][0] ;
 wire \line_cache[19][1] ;
 wire \line_cache[19][2] ;
 wire \line_cache[19][3] ;
 wire \line_cache[19][4] ;
 wire \line_cache[19][5] ;
 wire \line_cache[19][6] ;
 wire \line_cache[19][7] ;
 wire \line_cache[1][0] ;
 wire \line_cache[1][1] ;
 wire \line_cache[1][2] ;
 wire \line_cache[1][3] ;
 wire \line_cache[1][4] ;
 wire \line_cache[1][5] ;
 wire \line_cache[1][6] ;
 wire \line_cache[1][7] ;
 wire \line_cache[200][0] ;
 wire \line_cache[200][1] ;
 wire \line_cache[200][2] ;
 wire \line_cache[200][3] ;
 wire \line_cache[200][4] ;
 wire \line_cache[200][5] ;
 wire \line_cache[200][6] ;
 wire \line_cache[200][7] ;
 wire \line_cache[201][0] ;
 wire \line_cache[201][1] ;
 wire \line_cache[201][2] ;
 wire \line_cache[201][3] ;
 wire \line_cache[201][4] ;
 wire \line_cache[201][5] ;
 wire \line_cache[201][6] ;
 wire \line_cache[201][7] ;
 wire \line_cache[202][0] ;
 wire \line_cache[202][1] ;
 wire \line_cache[202][2] ;
 wire \line_cache[202][3] ;
 wire \line_cache[202][4] ;
 wire \line_cache[202][5] ;
 wire \line_cache[202][6] ;
 wire \line_cache[202][7] ;
 wire \line_cache[203][0] ;
 wire \line_cache[203][1] ;
 wire \line_cache[203][2] ;
 wire \line_cache[203][3] ;
 wire \line_cache[203][4] ;
 wire \line_cache[203][5] ;
 wire \line_cache[203][6] ;
 wire \line_cache[203][7] ;
 wire \line_cache[204][0] ;
 wire \line_cache[204][1] ;
 wire \line_cache[204][2] ;
 wire \line_cache[204][3] ;
 wire \line_cache[204][4] ;
 wire \line_cache[204][5] ;
 wire \line_cache[204][6] ;
 wire \line_cache[204][7] ;
 wire \line_cache[205][0] ;
 wire \line_cache[205][1] ;
 wire \line_cache[205][2] ;
 wire \line_cache[205][3] ;
 wire \line_cache[205][4] ;
 wire \line_cache[205][5] ;
 wire \line_cache[205][6] ;
 wire \line_cache[205][7] ;
 wire \line_cache[206][0] ;
 wire \line_cache[206][1] ;
 wire \line_cache[206][2] ;
 wire \line_cache[206][3] ;
 wire \line_cache[206][4] ;
 wire \line_cache[206][5] ;
 wire \line_cache[206][6] ;
 wire \line_cache[206][7] ;
 wire \line_cache[207][0] ;
 wire \line_cache[207][1] ;
 wire \line_cache[207][2] ;
 wire \line_cache[207][3] ;
 wire \line_cache[207][4] ;
 wire \line_cache[207][5] ;
 wire \line_cache[207][6] ;
 wire \line_cache[207][7] ;
 wire \line_cache[208][0] ;
 wire \line_cache[208][1] ;
 wire \line_cache[208][2] ;
 wire \line_cache[208][3] ;
 wire \line_cache[208][4] ;
 wire \line_cache[208][5] ;
 wire \line_cache[208][6] ;
 wire \line_cache[208][7] ;
 wire \line_cache[209][0] ;
 wire \line_cache[209][1] ;
 wire \line_cache[209][2] ;
 wire \line_cache[209][3] ;
 wire \line_cache[209][4] ;
 wire \line_cache[209][5] ;
 wire \line_cache[209][6] ;
 wire \line_cache[209][7] ;
 wire \line_cache[20][0] ;
 wire \line_cache[20][1] ;
 wire \line_cache[20][2] ;
 wire \line_cache[20][3] ;
 wire \line_cache[20][4] ;
 wire \line_cache[20][5] ;
 wire \line_cache[20][6] ;
 wire \line_cache[20][7] ;
 wire \line_cache[210][0] ;
 wire \line_cache[210][1] ;
 wire \line_cache[210][2] ;
 wire \line_cache[210][3] ;
 wire \line_cache[210][4] ;
 wire \line_cache[210][5] ;
 wire \line_cache[210][6] ;
 wire \line_cache[210][7] ;
 wire \line_cache[211][0] ;
 wire \line_cache[211][1] ;
 wire \line_cache[211][2] ;
 wire \line_cache[211][3] ;
 wire \line_cache[211][4] ;
 wire \line_cache[211][5] ;
 wire \line_cache[211][6] ;
 wire \line_cache[211][7] ;
 wire \line_cache[212][0] ;
 wire \line_cache[212][1] ;
 wire \line_cache[212][2] ;
 wire \line_cache[212][3] ;
 wire \line_cache[212][4] ;
 wire \line_cache[212][5] ;
 wire \line_cache[212][6] ;
 wire \line_cache[212][7] ;
 wire \line_cache[213][0] ;
 wire \line_cache[213][1] ;
 wire \line_cache[213][2] ;
 wire \line_cache[213][3] ;
 wire \line_cache[213][4] ;
 wire \line_cache[213][5] ;
 wire \line_cache[213][6] ;
 wire \line_cache[213][7] ;
 wire \line_cache[214][0] ;
 wire \line_cache[214][1] ;
 wire \line_cache[214][2] ;
 wire \line_cache[214][3] ;
 wire \line_cache[214][4] ;
 wire \line_cache[214][5] ;
 wire \line_cache[214][6] ;
 wire \line_cache[214][7] ;
 wire \line_cache[215][0] ;
 wire \line_cache[215][1] ;
 wire \line_cache[215][2] ;
 wire \line_cache[215][3] ;
 wire \line_cache[215][4] ;
 wire \line_cache[215][5] ;
 wire \line_cache[215][6] ;
 wire \line_cache[215][7] ;
 wire \line_cache[216][0] ;
 wire \line_cache[216][1] ;
 wire \line_cache[216][2] ;
 wire \line_cache[216][3] ;
 wire \line_cache[216][4] ;
 wire \line_cache[216][5] ;
 wire \line_cache[216][6] ;
 wire \line_cache[216][7] ;
 wire \line_cache[217][0] ;
 wire \line_cache[217][1] ;
 wire \line_cache[217][2] ;
 wire \line_cache[217][3] ;
 wire \line_cache[217][4] ;
 wire \line_cache[217][5] ;
 wire \line_cache[217][6] ;
 wire \line_cache[217][7] ;
 wire \line_cache[218][0] ;
 wire \line_cache[218][1] ;
 wire \line_cache[218][2] ;
 wire \line_cache[218][3] ;
 wire \line_cache[218][4] ;
 wire \line_cache[218][5] ;
 wire \line_cache[218][6] ;
 wire \line_cache[218][7] ;
 wire \line_cache[219][0] ;
 wire \line_cache[219][1] ;
 wire \line_cache[219][2] ;
 wire \line_cache[219][3] ;
 wire \line_cache[219][4] ;
 wire \line_cache[219][5] ;
 wire \line_cache[219][6] ;
 wire \line_cache[219][7] ;
 wire \line_cache[21][0] ;
 wire \line_cache[21][1] ;
 wire \line_cache[21][2] ;
 wire \line_cache[21][3] ;
 wire \line_cache[21][4] ;
 wire \line_cache[21][5] ;
 wire \line_cache[21][6] ;
 wire \line_cache[21][7] ;
 wire \line_cache[220][0] ;
 wire \line_cache[220][1] ;
 wire \line_cache[220][2] ;
 wire \line_cache[220][3] ;
 wire \line_cache[220][4] ;
 wire \line_cache[220][5] ;
 wire \line_cache[220][6] ;
 wire \line_cache[220][7] ;
 wire \line_cache[221][0] ;
 wire \line_cache[221][1] ;
 wire \line_cache[221][2] ;
 wire \line_cache[221][3] ;
 wire \line_cache[221][4] ;
 wire \line_cache[221][5] ;
 wire \line_cache[221][6] ;
 wire \line_cache[221][7] ;
 wire \line_cache[222][0] ;
 wire \line_cache[222][1] ;
 wire \line_cache[222][2] ;
 wire \line_cache[222][3] ;
 wire \line_cache[222][4] ;
 wire \line_cache[222][5] ;
 wire \line_cache[222][6] ;
 wire \line_cache[222][7] ;
 wire \line_cache[223][0] ;
 wire \line_cache[223][1] ;
 wire \line_cache[223][2] ;
 wire \line_cache[223][3] ;
 wire \line_cache[223][4] ;
 wire \line_cache[223][5] ;
 wire \line_cache[223][6] ;
 wire \line_cache[223][7] ;
 wire \line_cache[224][0] ;
 wire \line_cache[224][1] ;
 wire \line_cache[224][2] ;
 wire \line_cache[224][3] ;
 wire \line_cache[224][4] ;
 wire \line_cache[224][5] ;
 wire \line_cache[224][6] ;
 wire \line_cache[224][7] ;
 wire \line_cache[225][0] ;
 wire \line_cache[225][1] ;
 wire \line_cache[225][2] ;
 wire \line_cache[225][3] ;
 wire \line_cache[225][4] ;
 wire \line_cache[225][5] ;
 wire \line_cache[225][6] ;
 wire \line_cache[225][7] ;
 wire \line_cache[226][0] ;
 wire \line_cache[226][1] ;
 wire \line_cache[226][2] ;
 wire \line_cache[226][3] ;
 wire \line_cache[226][4] ;
 wire \line_cache[226][5] ;
 wire \line_cache[226][6] ;
 wire \line_cache[226][7] ;
 wire \line_cache[227][0] ;
 wire \line_cache[227][1] ;
 wire \line_cache[227][2] ;
 wire \line_cache[227][3] ;
 wire \line_cache[227][4] ;
 wire \line_cache[227][5] ;
 wire \line_cache[227][6] ;
 wire \line_cache[227][7] ;
 wire \line_cache[228][0] ;
 wire \line_cache[228][1] ;
 wire \line_cache[228][2] ;
 wire \line_cache[228][3] ;
 wire \line_cache[228][4] ;
 wire \line_cache[228][5] ;
 wire \line_cache[228][6] ;
 wire \line_cache[228][7] ;
 wire \line_cache[229][0] ;
 wire \line_cache[229][1] ;
 wire \line_cache[229][2] ;
 wire \line_cache[229][3] ;
 wire \line_cache[229][4] ;
 wire \line_cache[229][5] ;
 wire \line_cache[229][6] ;
 wire \line_cache[229][7] ;
 wire \line_cache[22][0] ;
 wire \line_cache[22][1] ;
 wire \line_cache[22][2] ;
 wire \line_cache[22][3] ;
 wire \line_cache[22][4] ;
 wire \line_cache[22][5] ;
 wire \line_cache[22][6] ;
 wire \line_cache[22][7] ;
 wire \line_cache[230][0] ;
 wire \line_cache[230][1] ;
 wire \line_cache[230][2] ;
 wire \line_cache[230][3] ;
 wire \line_cache[230][4] ;
 wire \line_cache[230][5] ;
 wire \line_cache[230][6] ;
 wire \line_cache[230][7] ;
 wire \line_cache[231][0] ;
 wire \line_cache[231][1] ;
 wire \line_cache[231][2] ;
 wire \line_cache[231][3] ;
 wire \line_cache[231][4] ;
 wire \line_cache[231][5] ;
 wire \line_cache[231][6] ;
 wire \line_cache[231][7] ;
 wire \line_cache[232][0] ;
 wire \line_cache[232][1] ;
 wire \line_cache[232][2] ;
 wire \line_cache[232][3] ;
 wire \line_cache[232][4] ;
 wire \line_cache[232][5] ;
 wire \line_cache[232][6] ;
 wire \line_cache[232][7] ;
 wire \line_cache[233][0] ;
 wire \line_cache[233][1] ;
 wire \line_cache[233][2] ;
 wire \line_cache[233][3] ;
 wire \line_cache[233][4] ;
 wire \line_cache[233][5] ;
 wire \line_cache[233][6] ;
 wire \line_cache[233][7] ;
 wire \line_cache[234][0] ;
 wire \line_cache[234][1] ;
 wire \line_cache[234][2] ;
 wire \line_cache[234][3] ;
 wire \line_cache[234][4] ;
 wire \line_cache[234][5] ;
 wire \line_cache[234][6] ;
 wire \line_cache[234][7] ;
 wire \line_cache[235][0] ;
 wire \line_cache[235][1] ;
 wire \line_cache[235][2] ;
 wire \line_cache[235][3] ;
 wire \line_cache[235][4] ;
 wire \line_cache[235][5] ;
 wire \line_cache[235][6] ;
 wire \line_cache[235][7] ;
 wire \line_cache[236][0] ;
 wire \line_cache[236][1] ;
 wire \line_cache[236][2] ;
 wire \line_cache[236][3] ;
 wire \line_cache[236][4] ;
 wire \line_cache[236][5] ;
 wire \line_cache[236][6] ;
 wire \line_cache[236][7] ;
 wire \line_cache[237][0] ;
 wire \line_cache[237][1] ;
 wire \line_cache[237][2] ;
 wire \line_cache[237][3] ;
 wire \line_cache[237][4] ;
 wire \line_cache[237][5] ;
 wire \line_cache[237][6] ;
 wire \line_cache[237][7] ;
 wire \line_cache[238][0] ;
 wire \line_cache[238][1] ;
 wire \line_cache[238][2] ;
 wire \line_cache[238][3] ;
 wire \line_cache[238][4] ;
 wire \line_cache[238][5] ;
 wire \line_cache[238][6] ;
 wire \line_cache[238][7] ;
 wire \line_cache[239][0] ;
 wire \line_cache[239][1] ;
 wire \line_cache[239][2] ;
 wire \line_cache[239][3] ;
 wire \line_cache[239][4] ;
 wire \line_cache[239][5] ;
 wire \line_cache[239][6] ;
 wire \line_cache[239][7] ;
 wire \line_cache[23][0] ;
 wire \line_cache[23][1] ;
 wire \line_cache[23][2] ;
 wire \line_cache[23][3] ;
 wire \line_cache[23][4] ;
 wire \line_cache[23][5] ;
 wire \line_cache[23][6] ;
 wire \line_cache[23][7] ;
 wire \line_cache[240][0] ;
 wire \line_cache[240][1] ;
 wire \line_cache[240][2] ;
 wire \line_cache[240][3] ;
 wire \line_cache[240][4] ;
 wire \line_cache[240][5] ;
 wire \line_cache[240][6] ;
 wire \line_cache[240][7] ;
 wire \line_cache[241][0] ;
 wire \line_cache[241][1] ;
 wire \line_cache[241][2] ;
 wire \line_cache[241][3] ;
 wire \line_cache[241][4] ;
 wire \line_cache[241][5] ;
 wire \line_cache[241][6] ;
 wire \line_cache[241][7] ;
 wire \line_cache[242][0] ;
 wire \line_cache[242][1] ;
 wire \line_cache[242][2] ;
 wire \line_cache[242][3] ;
 wire \line_cache[242][4] ;
 wire \line_cache[242][5] ;
 wire \line_cache[242][6] ;
 wire \line_cache[242][7] ;
 wire \line_cache[243][0] ;
 wire \line_cache[243][1] ;
 wire \line_cache[243][2] ;
 wire \line_cache[243][3] ;
 wire \line_cache[243][4] ;
 wire \line_cache[243][5] ;
 wire \line_cache[243][6] ;
 wire \line_cache[243][7] ;
 wire \line_cache[244][0] ;
 wire \line_cache[244][1] ;
 wire \line_cache[244][2] ;
 wire \line_cache[244][3] ;
 wire \line_cache[244][4] ;
 wire \line_cache[244][5] ;
 wire \line_cache[244][6] ;
 wire \line_cache[244][7] ;
 wire \line_cache[245][0] ;
 wire \line_cache[245][1] ;
 wire \line_cache[245][2] ;
 wire \line_cache[245][3] ;
 wire \line_cache[245][4] ;
 wire \line_cache[245][5] ;
 wire \line_cache[245][6] ;
 wire \line_cache[245][7] ;
 wire \line_cache[246][0] ;
 wire \line_cache[246][1] ;
 wire \line_cache[246][2] ;
 wire \line_cache[246][3] ;
 wire \line_cache[246][4] ;
 wire \line_cache[246][5] ;
 wire \line_cache[246][6] ;
 wire \line_cache[246][7] ;
 wire \line_cache[247][0] ;
 wire \line_cache[247][1] ;
 wire \line_cache[247][2] ;
 wire \line_cache[247][3] ;
 wire \line_cache[247][4] ;
 wire \line_cache[247][5] ;
 wire \line_cache[247][6] ;
 wire \line_cache[247][7] ;
 wire \line_cache[248][0] ;
 wire \line_cache[248][1] ;
 wire \line_cache[248][2] ;
 wire \line_cache[248][3] ;
 wire \line_cache[248][4] ;
 wire \line_cache[248][5] ;
 wire \line_cache[248][6] ;
 wire \line_cache[248][7] ;
 wire \line_cache[249][0] ;
 wire \line_cache[249][1] ;
 wire \line_cache[249][2] ;
 wire \line_cache[249][3] ;
 wire \line_cache[249][4] ;
 wire \line_cache[249][5] ;
 wire \line_cache[249][6] ;
 wire \line_cache[249][7] ;
 wire \line_cache[24][0] ;
 wire \line_cache[24][1] ;
 wire \line_cache[24][2] ;
 wire \line_cache[24][3] ;
 wire \line_cache[24][4] ;
 wire \line_cache[24][5] ;
 wire \line_cache[24][6] ;
 wire \line_cache[24][7] ;
 wire \line_cache[250][0] ;
 wire \line_cache[250][1] ;
 wire \line_cache[250][2] ;
 wire \line_cache[250][3] ;
 wire \line_cache[250][4] ;
 wire \line_cache[250][5] ;
 wire \line_cache[250][6] ;
 wire \line_cache[250][7] ;
 wire \line_cache[251][0] ;
 wire \line_cache[251][1] ;
 wire \line_cache[251][2] ;
 wire \line_cache[251][3] ;
 wire \line_cache[251][4] ;
 wire \line_cache[251][5] ;
 wire \line_cache[251][6] ;
 wire \line_cache[251][7] ;
 wire \line_cache[252][0] ;
 wire \line_cache[252][1] ;
 wire \line_cache[252][2] ;
 wire \line_cache[252][3] ;
 wire \line_cache[252][4] ;
 wire \line_cache[252][5] ;
 wire \line_cache[252][6] ;
 wire \line_cache[252][7] ;
 wire \line_cache[253][0] ;
 wire \line_cache[253][1] ;
 wire \line_cache[253][2] ;
 wire \line_cache[253][3] ;
 wire \line_cache[253][4] ;
 wire \line_cache[253][5] ;
 wire \line_cache[253][6] ;
 wire \line_cache[253][7] ;
 wire \line_cache[254][0] ;
 wire \line_cache[254][1] ;
 wire \line_cache[254][2] ;
 wire \line_cache[254][3] ;
 wire \line_cache[254][4] ;
 wire \line_cache[254][5] ;
 wire \line_cache[254][6] ;
 wire \line_cache[254][7] ;
 wire \line_cache[255][0] ;
 wire \line_cache[255][1] ;
 wire \line_cache[255][2] ;
 wire \line_cache[255][3] ;
 wire \line_cache[255][4] ;
 wire \line_cache[255][5] ;
 wire \line_cache[255][6] ;
 wire \line_cache[255][7] ;
 wire \line_cache[256][0] ;
 wire \line_cache[256][1] ;
 wire \line_cache[256][2] ;
 wire \line_cache[256][3] ;
 wire \line_cache[256][4] ;
 wire \line_cache[256][5] ;
 wire \line_cache[256][6] ;
 wire \line_cache[256][7] ;
 wire \line_cache[257][0] ;
 wire \line_cache[257][1] ;
 wire \line_cache[257][2] ;
 wire \line_cache[257][3] ;
 wire \line_cache[257][4] ;
 wire \line_cache[257][5] ;
 wire \line_cache[257][6] ;
 wire \line_cache[257][7] ;
 wire \line_cache[258][0] ;
 wire \line_cache[258][1] ;
 wire \line_cache[258][2] ;
 wire \line_cache[258][3] ;
 wire \line_cache[258][4] ;
 wire \line_cache[258][5] ;
 wire \line_cache[258][6] ;
 wire \line_cache[258][7] ;
 wire \line_cache[259][0] ;
 wire \line_cache[259][1] ;
 wire \line_cache[259][2] ;
 wire \line_cache[259][3] ;
 wire \line_cache[259][4] ;
 wire \line_cache[259][5] ;
 wire \line_cache[259][6] ;
 wire \line_cache[259][7] ;
 wire \line_cache[25][0] ;
 wire \line_cache[25][1] ;
 wire \line_cache[25][2] ;
 wire \line_cache[25][3] ;
 wire \line_cache[25][4] ;
 wire \line_cache[25][5] ;
 wire \line_cache[25][6] ;
 wire \line_cache[25][7] ;
 wire \line_cache[260][0] ;
 wire \line_cache[260][1] ;
 wire \line_cache[260][2] ;
 wire \line_cache[260][3] ;
 wire \line_cache[260][4] ;
 wire \line_cache[260][5] ;
 wire \line_cache[260][6] ;
 wire \line_cache[260][7] ;
 wire \line_cache[261][0] ;
 wire \line_cache[261][1] ;
 wire \line_cache[261][2] ;
 wire \line_cache[261][3] ;
 wire \line_cache[261][4] ;
 wire \line_cache[261][5] ;
 wire \line_cache[261][6] ;
 wire \line_cache[261][7] ;
 wire \line_cache[262][0] ;
 wire \line_cache[262][1] ;
 wire \line_cache[262][2] ;
 wire \line_cache[262][3] ;
 wire \line_cache[262][4] ;
 wire \line_cache[262][5] ;
 wire \line_cache[262][6] ;
 wire \line_cache[262][7] ;
 wire \line_cache[263][0] ;
 wire \line_cache[263][1] ;
 wire \line_cache[263][2] ;
 wire \line_cache[263][3] ;
 wire \line_cache[263][4] ;
 wire \line_cache[263][5] ;
 wire \line_cache[263][6] ;
 wire \line_cache[263][7] ;
 wire \line_cache[264][0] ;
 wire \line_cache[264][1] ;
 wire \line_cache[264][2] ;
 wire \line_cache[264][3] ;
 wire \line_cache[264][4] ;
 wire \line_cache[264][5] ;
 wire \line_cache[264][6] ;
 wire \line_cache[264][7] ;
 wire \line_cache[265][0] ;
 wire \line_cache[265][1] ;
 wire \line_cache[265][2] ;
 wire \line_cache[265][3] ;
 wire \line_cache[265][4] ;
 wire \line_cache[265][5] ;
 wire \line_cache[265][6] ;
 wire \line_cache[265][7] ;
 wire \line_cache[266][0] ;
 wire \line_cache[266][1] ;
 wire \line_cache[266][2] ;
 wire \line_cache[266][3] ;
 wire \line_cache[266][4] ;
 wire \line_cache[266][5] ;
 wire \line_cache[266][6] ;
 wire \line_cache[266][7] ;
 wire \line_cache[267][0] ;
 wire \line_cache[267][1] ;
 wire \line_cache[267][2] ;
 wire \line_cache[267][3] ;
 wire \line_cache[267][4] ;
 wire \line_cache[267][5] ;
 wire \line_cache[267][6] ;
 wire \line_cache[267][7] ;
 wire \line_cache[268][0] ;
 wire \line_cache[268][1] ;
 wire \line_cache[268][2] ;
 wire \line_cache[268][3] ;
 wire \line_cache[268][4] ;
 wire \line_cache[268][5] ;
 wire \line_cache[268][6] ;
 wire \line_cache[268][7] ;
 wire \line_cache[269][0] ;
 wire \line_cache[269][1] ;
 wire \line_cache[269][2] ;
 wire \line_cache[269][3] ;
 wire \line_cache[269][4] ;
 wire \line_cache[269][5] ;
 wire \line_cache[269][6] ;
 wire \line_cache[269][7] ;
 wire \line_cache[26][0] ;
 wire \line_cache[26][1] ;
 wire \line_cache[26][2] ;
 wire \line_cache[26][3] ;
 wire \line_cache[26][4] ;
 wire \line_cache[26][5] ;
 wire \line_cache[26][6] ;
 wire \line_cache[26][7] ;
 wire \line_cache[270][0] ;
 wire \line_cache[270][1] ;
 wire \line_cache[270][2] ;
 wire \line_cache[270][3] ;
 wire \line_cache[270][4] ;
 wire \line_cache[270][5] ;
 wire \line_cache[270][6] ;
 wire \line_cache[270][7] ;
 wire \line_cache[271][0] ;
 wire \line_cache[271][1] ;
 wire \line_cache[271][2] ;
 wire \line_cache[271][3] ;
 wire \line_cache[271][4] ;
 wire \line_cache[271][5] ;
 wire \line_cache[271][6] ;
 wire \line_cache[271][7] ;
 wire \line_cache[272][0] ;
 wire \line_cache[272][1] ;
 wire \line_cache[272][2] ;
 wire \line_cache[272][3] ;
 wire \line_cache[272][4] ;
 wire \line_cache[272][5] ;
 wire \line_cache[272][6] ;
 wire \line_cache[272][7] ;
 wire \line_cache[273][0] ;
 wire \line_cache[273][1] ;
 wire \line_cache[273][2] ;
 wire \line_cache[273][3] ;
 wire \line_cache[273][4] ;
 wire \line_cache[273][5] ;
 wire \line_cache[273][6] ;
 wire \line_cache[273][7] ;
 wire \line_cache[274][0] ;
 wire \line_cache[274][1] ;
 wire \line_cache[274][2] ;
 wire \line_cache[274][3] ;
 wire \line_cache[274][4] ;
 wire \line_cache[274][5] ;
 wire \line_cache[274][6] ;
 wire \line_cache[274][7] ;
 wire \line_cache[275][0] ;
 wire \line_cache[275][1] ;
 wire \line_cache[275][2] ;
 wire \line_cache[275][3] ;
 wire \line_cache[275][4] ;
 wire \line_cache[275][5] ;
 wire \line_cache[275][6] ;
 wire \line_cache[275][7] ;
 wire \line_cache[276][0] ;
 wire \line_cache[276][1] ;
 wire \line_cache[276][2] ;
 wire \line_cache[276][3] ;
 wire \line_cache[276][4] ;
 wire \line_cache[276][5] ;
 wire \line_cache[276][6] ;
 wire \line_cache[276][7] ;
 wire \line_cache[277][0] ;
 wire \line_cache[277][1] ;
 wire \line_cache[277][2] ;
 wire \line_cache[277][3] ;
 wire \line_cache[277][4] ;
 wire \line_cache[277][5] ;
 wire \line_cache[277][6] ;
 wire \line_cache[277][7] ;
 wire \line_cache[278][0] ;
 wire \line_cache[278][1] ;
 wire \line_cache[278][2] ;
 wire \line_cache[278][3] ;
 wire \line_cache[278][4] ;
 wire \line_cache[278][5] ;
 wire \line_cache[278][6] ;
 wire \line_cache[278][7] ;
 wire \line_cache[279][0] ;
 wire \line_cache[279][1] ;
 wire \line_cache[279][2] ;
 wire \line_cache[279][3] ;
 wire \line_cache[279][4] ;
 wire \line_cache[279][5] ;
 wire \line_cache[279][6] ;
 wire \line_cache[279][7] ;
 wire \line_cache[27][0] ;
 wire \line_cache[27][1] ;
 wire \line_cache[27][2] ;
 wire \line_cache[27][3] ;
 wire \line_cache[27][4] ;
 wire \line_cache[27][5] ;
 wire \line_cache[27][6] ;
 wire \line_cache[27][7] ;
 wire \line_cache[280][0] ;
 wire \line_cache[280][1] ;
 wire \line_cache[280][2] ;
 wire \line_cache[280][3] ;
 wire \line_cache[280][4] ;
 wire \line_cache[280][5] ;
 wire \line_cache[280][6] ;
 wire \line_cache[280][7] ;
 wire \line_cache[281][0] ;
 wire \line_cache[281][1] ;
 wire \line_cache[281][2] ;
 wire \line_cache[281][3] ;
 wire \line_cache[281][4] ;
 wire \line_cache[281][5] ;
 wire \line_cache[281][6] ;
 wire \line_cache[281][7] ;
 wire \line_cache[282][0] ;
 wire \line_cache[282][1] ;
 wire \line_cache[282][2] ;
 wire \line_cache[282][3] ;
 wire \line_cache[282][4] ;
 wire \line_cache[282][5] ;
 wire \line_cache[282][6] ;
 wire \line_cache[282][7] ;
 wire \line_cache[283][0] ;
 wire \line_cache[283][1] ;
 wire \line_cache[283][2] ;
 wire \line_cache[283][3] ;
 wire \line_cache[283][4] ;
 wire \line_cache[283][5] ;
 wire \line_cache[283][6] ;
 wire \line_cache[283][7] ;
 wire \line_cache[284][0] ;
 wire \line_cache[284][1] ;
 wire \line_cache[284][2] ;
 wire \line_cache[284][3] ;
 wire \line_cache[284][4] ;
 wire \line_cache[284][5] ;
 wire \line_cache[284][6] ;
 wire \line_cache[284][7] ;
 wire \line_cache[285][0] ;
 wire \line_cache[285][1] ;
 wire \line_cache[285][2] ;
 wire \line_cache[285][3] ;
 wire \line_cache[285][4] ;
 wire \line_cache[285][5] ;
 wire \line_cache[285][6] ;
 wire \line_cache[285][7] ;
 wire \line_cache[286][0] ;
 wire \line_cache[286][1] ;
 wire \line_cache[286][2] ;
 wire \line_cache[286][3] ;
 wire \line_cache[286][4] ;
 wire \line_cache[286][5] ;
 wire \line_cache[286][6] ;
 wire \line_cache[286][7] ;
 wire \line_cache[287][0] ;
 wire \line_cache[287][1] ;
 wire \line_cache[287][2] ;
 wire \line_cache[287][3] ;
 wire \line_cache[287][4] ;
 wire \line_cache[287][5] ;
 wire \line_cache[287][6] ;
 wire \line_cache[287][7] ;
 wire \line_cache[288][0] ;
 wire \line_cache[288][1] ;
 wire \line_cache[288][2] ;
 wire \line_cache[288][3] ;
 wire \line_cache[288][4] ;
 wire \line_cache[288][5] ;
 wire \line_cache[288][6] ;
 wire \line_cache[288][7] ;
 wire \line_cache[289][0] ;
 wire \line_cache[289][1] ;
 wire \line_cache[289][2] ;
 wire \line_cache[289][3] ;
 wire \line_cache[289][4] ;
 wire \line_cache[289][5] ;
 wire \line_cache[289][6] ;
 wire \line_cache[289][7] ;
 wire \line_cache[28][0] ;
 wire \line_cache[28][1] ;
 wire \line_cache[28][2] ;
 wire \line_cache[28][3] ;
 wire \line_cache[28][4] ;
 wire \line_cache[28][5] ;
 wire \line_cache[28][6] ;
 wire \line_cache[28][7] ;
 wire \line_cache[290][0] ;
 wire \line_cache[290][1] ;
 wire \line_cache[290][2] ;
 wire \line_cache[290][3] ;
 wire \line_cache[290][4] ;
 wire \line_cache[290][5] ;
 wire \line_cache[290][6] ;
 wire \line_cache[290][7] ;
 wire \line_cache[291][0] ;
 wire \line_cache[291][1] ;
 wire \line_cache[291][2] ;
 wire \line_cache[291][3] ;
 wire \line_cache[291][4] ;
 wire \line_cache[291][5] ;
 wire \line_cache[291][6] ;
 wire \line_cache[291][7] ;
 wire \line_cache[292][0] ;
 wire \line_cache[292][1] ;
 wire \line_cache[292][2] ;
 wire \line_cache[292][3] ;
 wire \line_cache[292][4] ;
 wire \line_cache[292][5] ;
 wire \line_cache[292][6] ;
 wire \line_cache[292][7] ;
 wire \line_cache[293][0] ;
 wire \line_cache[293][1] ;
 wire \line_cache[293][2] ;
 wire \line_cache[293][3] ;
 wire \line_cache[293][4] ;
 wire \line_cache[293][5] ;
 wire \line_cache[293][6] ;
 wire \line_cache[293][7] ;
 wire \line_cache[294][0] ;
 wire \line_cache[294][1] ;
 wire \line_cache[294][2] ;
 wire \line_cache[294][3] ;
 wire \line_cache[294][4] ;
 wire \line_cache[294][5] ;
 wire \line_cache[294][6] ;
 wire \line_cache[294][7] ;
 wire \line_cache[295][0] ;
 wire \line_cache[295][1] ;
 wire \line_cache[295][2] ;
 wire \line_cache[295][3] ;
 wire \line_cache[295][4] ;
 wire \line_cache[295][5] ;
 wire \line_cache[295][6] ;
 wire \line_cache[295][7] ;
 wire \line_cache[296][0] ;
 wire \line_cache[296][1] ;
 wire \line_cache[296][2] ;
 wire \line_cache[296][3] ;
 wire \line_cache[296][4] ;
 wire \line_cache[296][5] ;
 wire \line_cache[296][6] ;
 wire \line_cache[296][7] ;
 wire \line_cache[297][0] ;
 wire \line_cache[297][1] ;
 wire \line_cache[297][2] ;
 wire \line_cache[297][3] ;
 wire \line_cache[297][4] ;
 wire \line_cache[297][5] ;
 wire \line_cache[297][6] ;
 wire \line_cache[297][7] ;
 wire \line_cache[298][0] ;
 wire \line_cache[298][1] ;
 wire \line_cache[298][2] ;
 wire \line_cache[298][3] ;
 wire \line_cache[298][4] ;
 wire \line_cache[298][5] ;
 wire \line_cache[298][6] ;
 wire \line_cache[298][7] ;
 wire \line_cache[299][0] ;
 wire \line_cache[299][1] ;
 wire \line_cache[299][2] ;
 wire \line_cache[299][3] ;
 wire \line_cache[299][4] ;
 wire \line_cache[299][5] ;
 wire \line_cache[299][6] ;
 wire \line_cache[299][7] ;
 wire \line_cache[29][0] ;
 wire \line_cache[29][1] ;
 wire \line_cache[29][2] ;
 wire \line_cache[29][3] ;
 wire \line_cache[29][4] ;
 wire \line_cache[29][5] ;
 wire \line_cache[29][6] ;
 wire \line_cache[29][7] ;
 wire \line_cache[2][0] ;
 wire \line_cache[2][1] ;
 wire \line_cache[2][2] ;
 wire \line_cache[2][3] ;
 wire \line_cache[2][4] ;
 wire \line_cache[2][5] ;
 wire \line_cache[2][6] ;
 wire \line_cache[2][7] ;
 wire \line_cache[300][0] ;
 wire \line_cache[300][1] ;
 wire \line_cache[300][2] ;
 wire \line_cache[300][3] ;
 wire \line_cache[300][4] ;
 wire \line_cache[300][5] ;
 wire \line_cache[300][6] ;
 wire \line_cache[300][7] ;
 wire \line_cache[301][0] ;
 wire \line_cache[301][1] ;
 wire \line_cache[301][2] ;
 wire \line_cache[301][3] ;
 wire \line_cache[301][4] ;
 wire \line_cache[301][5] ;
 wire \line_cache[301][6] ;
 wire \line_cache[301][7] ;
 wire \line_cache[302][0] ;
 wire \line_cache[302][1] ;
 wire \line_cache[302][2] ;
 wire \line_cache[302][3] ;
 wire \line_cache[302][4] ;
 wire \line_cache[302][5] ;
 wire \line_cache[302][6] ;
 wire \line_cache[302][7] ;
 wire \line_cache[303][0] ;
 wire \line_cache[303][1] ;
 wire \line_cache[303][2] ;
 wire \line_cache[303][3] ;
 wire \line_cache[303][4] ;
 wire \line_cache[303][5] ;
 wire \line_cache[303][6] ;
 wire \line_cache[303][7] ;
 wire \line_cache[304][0] ;
 wire \line_cache[304][1] ;
 wire \line_cache[304][2] ;
 wire \line_cache[304][3] ;
 wire \line_cache[304][4] ;
 wire \line_cache[304][5] ;
 wire \line_cache[304][6] ;
 wire \line_cache[304][7] ;
 wire \line_cache[305][0] ;
 wire \line_cache[305][1] ;
 wire \line_cache[305][2] ;
 wire \line_cache[305][3] ;
 wire \line_cache[305][4] ;
 wire \line_cache[305][5] ;
 wire \line_cache[305][6] ;
 wire \line_cache[305][7] ;
 wire \line_cache[306][0] ;
 wire \line_cache[306][1] ;
 wire \line_cache[306][2] ;
 wire \line_cache[306][3] ;
 wire \line_cache[306][4] ;
 wire \line_cache[306][5] ;
 wire \line_cache[306][6] ;
 wire \line_cache[306][7] ;
 wire \line_cache[307][0] ;
 wire \line_cache[307][1] ;
 wire \line_cache[307][2] ;
 wire \line_cache[307][3] ;
 wire \line_cache[307][4] ;
 wire \line_cache[307][5] ;
 wire \line_cache[307][6] ;
 wire \line_cache[307][7] ;
 wire \line_cache[308][0] ;
 wire \line_cache[308][1] ;
 wire \line_cache[308][2] ;
 wire \line_cache[308][3] ;
 wire \line_cache[308][4] ;
 wire \line_cache[308][5] ;
 wire \line_cache[308][6] ;
 wire \line_cache[308][7] ;
 wire \line_cache[309][0] ;
 wire \line_cache[309][1] ;
 wire \line_cache[309][2] ;
 wire \line_cache[309][3] ;
 wire \line_cache[309][4] ;
 wire \line_cache[309][5] ;
 wire \line_cache[309][6] ;
 wire \line_cache[309][7] ;
 wire \line_cache[30][0] ;
 wire \line_cache[30][1] ;
 wire \line_cache[30][2] ;
 wire \line_cache[30][3] ;
 wire \line_cache[30][4] ;
 wire \line_cache[30][5] ;
 wire \line_cache[30][6] ;
 wire \line_cache[30][7] ;
 wire \line_cache[310][0] ;
 wire \line_cache[310][1] ;
 wire \line_cache[310][2] ;
 wire \line_cache[310][3] ;
 wire \line_cache[310][4] ;
 wire \line_cache[310][5] ;
 wire \line_cache[310][6] ;
 wire \line_cache[310][7] ;
 wire \line_cache[311][0] ;
 wire \line_cache[311][1] ;
 wire \line_cache[311][2] ;
 wire \line_cache[311][3] ;
 wire \line_cache[311][4] ;
 wire \line_cache[311][5] ;
 wire \line_cache[311][6] ;
 wire \line_cache[311][7] ;
 wire \line_cache[312][0] ;
 wire \line_cache[312][1] ;
 wire \line_cache[312][2] ;
 wire \line_cache[312][3] ;
 wire \line_cache[312][4] ;
 wire \line_cache[312][5] ;
 wire \line_cache[312][6] ;
 wire \line_cache[312][7] ;
 wire \line_cache[313][0] ;
 wire \line_cache[313][1] ;
 wire \line_cache[313][2] ;
 wire \line_cache[313][3] ;
 wire \line_cache[313][4] ;
 wire \line_cache[313][5] ;
 wire \line_cache[313][6] ;
 wire \line_cache[313][7] ;
 wire \line_cache[314][0] ;
 wire \line_cache[314][1] ;
 wire \line_cache[314][2] ;
 wire \line_cache[314][3] ;
 wire \line_cache[314][4] ;
 wire \line_cache[314][5] ;
 wire \line_cache[314][6] ;
 wire \line_cache[314][7] ;
 wire \line_cache[315][0] ;
 wire \line_cache[315][1] ;
 wire \line_cache[315][2] ;
 wire \line_cache[315][3] ;
 wire \line_cache[315][4] ;
 wire \line_cache[315][5] ;
 wire \line_cache[315][6] ;
 wire \line_cache[315][7] ;
 wire \line_cache[316][0] ;
 wire \line_cache[316][1] ;
 wire \line_cache[316][2] ;
 wire \line_cache[316][3] ;
 wire \line_cache[316][4] ;
 wire \line_cache[316][5] ;
 wire \line_cache[316][6] ;
 wire \line_cache[316][7] ;
 wire \line_cache[317][0] ;
 wire \line_cache[317][1] ;
 wire \line_cache[317][2] ;
 wire \line_cache[317][3] ;
 wire \line_cache[317][4] ;
 wire \line_cache[317][5] ;
 wire \line_cache[317][6] ;
 wire \line_cache[317][7] ;
 wire \line_cache[318][0] ;
 wire \line_cache[318][1] ;
 wire \line_cache[318][2] ;
 wire \line_cache[318][3] ;
 wire \line_cache[318][4] ;
 wire \line_cache[318][5] ;
 wire \line_cache[318][6] ;
 wire \line_cache[318][7] ;
 wire \line_cache[319][0] ;
 wire \line_cache[319][1] ;
 wire \line_cache[319][2] ;
 wire \line_cache[319][3] ;
 wire \line_cache[319][4] ;
 wire \line_cache[319][5] ;
 wire \line_cache[319][6] ;
 wire \line_cache[319][7] ;
 wire \line_cache[31][0] ;
 wire \line_cache[31][1] ;
 wire \line_cache[31][2] ;
 wire \line_cache[31][3] ;
 wire \line_cache[31][4] ;
 wire \line_cache[31][5] ;
 wire \line_cache[31][6] ;
 wire \line_cache[31][7] ;
 wire \line_cache[32][0] ;
 wire \line_cache[32][1] ;
 wire \line_cache[32][2] ;
 wire \line_cache[32][3] ;
 wire \line_cache[32][4] ;
 wire \line_cache[32][5] ;
 wire \line_cache[32][6] ;
 wire \line_cache[32][7] ;
 wire \line_cache[33][0] ;
 wire \line_cache[33][1] ;
 wire \line_cache[33][2] ;
 wire \line_cache[33][3] ;
 wire \line_cache[33][4] ;
 wire \line_cache[33][5] ;
 wire \line_cache[33][6] ;
 wire \line_cache[33][7] ;
 wire \line_cache[34][0] ;
 wire \line_cache[34][1] ;
 wire \line_cache[34][2] ;
 wire \line_cache[34][3] ;
 wire \line_cache[34][4] ;
 wire \line_cache[34][5] ;
 wire \line_cache[34][6] ;
 wire \line_cache[34][7] ;
 wire \line_cache[35][0] ;
 wire \line_cache[35][1] ;
 wire \line_cache[35][2] ;
 wire \line_cache[35][3] ;
 wire \line_cache[35][4] ;
 wire \line_cache[35][5] ;
 wire \line_cache[35][6] ;
 wire \line_cache[35][7] ;
 wire \line_cache[36][0] ;
 wire \line_cache[36][1] ;
 wire \line_cache[36][2] ;
 wire \line_cache[36][3] ;
 wire \line_cache[36][4] ;
 wire \line_cache[36][5] ;
 wire \line_cache[36][6] ;
 wire \line_cache[36][7] ;
 wire \line_cache[37][0] ;
 wire \line_cache[37][1] ;
 wire \line_cache[37][2] ;
 wire \line_cache[37][3] ;
 wire \line_cache[37][4] ;
 wire \line_cache[37][5] ;
 wire \line_cache[37][6] ;
 wire \line_cache[37][7] ;
 wire \line_cache[38][0] ;
 wire \line_cache[38][1] ;
 wire \line_cache[38][2] ;
 wire \line_cache[38][3] ;
 wire \line_cache[38][4] ;
 wire \line_cache[38][5] ;
 wire \line_cache[38][6] ;
 wire \line_cache[38][7] ;
 wire \line_cache[39][0] ;
 wire \line_cache[39][1] ;
 wire \line_cache[39][2] ;
 wire \line_cache[39][3] ;
 wire \line_cache[39][4] ;
 wire \line_cache[39][5] ;
 wire \line_cache[39][6] ;
 wire \line_cache[39][7] ;
 wire \line_cache[3][0] ;
 wire \line_cache[3][1] ;
 wire \line_cache[3][2] ;
 wire \line_cache[3][3] ;
 wire \line_cache[3][4] ;
 wire \line_cache[3][5] ;
 wire \line_cache[3][6] ;
 wire \line_cache[3][7] ;
 wire \line_cache[40][0] ;
 wire \line_cache[40][1] ;
 wire \line_cache[40][2] ;
 wire \line_cache[40][3] ;
 wire \line_cache[40][4] ;
 wire \line_cache[40][5] ;
 wire \line_cache[40][6] ;
 wire \line_cache[40][7] ;
 wire \line_cache[41][0] ;
 wire \line_cache[41][1] ;
 wire \line_cache[41][2] ;
 wire \line_cache[41][3] ;
 wire \line_cache[41][4] ;
 wire \line_cache[41][5] ;
 wire \line_cache[41][6] ;
 wire \line_cache[41][7] ;
 wire \line_cache[42][0] ;
 wire \line_cache[42][1] ;
 wire \line_cache[42][2] ;
 wire \line_cache[42][3] ;
 wire \line_cache[42][4] ;
 wire \line_cache[42][5] ;
 wire \line_cache[42][6] ;
 wire \line_cache[42][7] ;
 wire \line_cache[43][0] ;
 wire \line_cache[43][1] ;
 wire \line_cache[43][2] ;
 wire \line_cache[43][3] ;
 wire \line_cache[43][4] ;
 wire \line_cache[43][5] ;
 wire \line_cache[43][6] ;
 wire \line_cache[43][7] ;
 wire \line_cache[44][0] ;
 wire \line_cache[44][1] ;
 wire \line_cache[44][2] ;
 wire \line_cache[44][3] ;
 wire \line_cache[44][4] ;
 wire \line_cache[44][5] ;
 wire \line_cache[44][6] ;
 wire \line_cache[44][7] ;
 wire \line_cache[45][0] ;
 wire \line_cache[45][1] ;
 wire \line_cache[45][2] ;
 wire \line_cache[45][3] ;
 wire \line_cache[45][4] ;
 wire \line_cache[45][5] ;
 wire \line_cache[45][6] ;
 wire \line_cache[45][7] ;
 wire \line_cache[46][0] ;
 wire \line_cache[46][1] ;
 wire \line_cache[46][2] ;
 wire \line_cache[46][3] ;
 wire \line_cache[46][4] ;
 wire \line_cache[46][5] ;
 wire \line_cache[46][6] ;
 wire \line_cache[46][7] ;
 wire \line_cache[47][0] ;
 wire \line_cache[47][1] ;
 wire \line_cache[47][2] ;
 wire \line_cache[47][3] ;
 wire \line_cache[47][4] ;
 wire \line_cache[47][5] ;
 wire \line_cache[47][6] ;
 wire \line_cache[47][7] ;
 wire \line_cache[48][0] ;
 wire \line_cache[48][1] ;
 wire \line_cache[48][2] ;
 wire \line_cache[48][3] ;
 wire \line_cache[48][4] ;
 wire \line_cache[48][5] ;
 wire \line_cache[48][6] ;
 wire \line_cache[48][7] ;
 wire \line_cache[49][0] ;
 wire \line_cache[49][1] ;
 wire \line_cache[49][2] ;
 wire \line_cache[49][3] ;
 wire \line_cache[49][4] ;
 wire \line_cache[49][5] ;
 wire \line_cache[49][6] ;
 wire \line_cache[49][7] ;
 wire \line_cache[4][0] ;
 wire \line_cache[4][1] ;
 wire \line_cache[4][2] ;
 wire \line_cache[4][3] ;
 wire \line_cache[4][4] ;
 wire \line_cache[4][5] ;
 wire \line_cache[4][6] ;
 wire \line_cache[4][7] ;
 wire \line_cache[50][0] ;
 wire \line_cache[50][1] ;
 wire \line_cache[50][2] ;
 wire \line_cache[50][3] ;
 wire \line_cache[50][4] ;
 wire \line_cache[50][5] ;
 wire \line_cache[50][6] ;
 wire \line_cache[50][7] ;
 wire \line_cache[51][0] ;
 wire \line_cache[51][1] ;
 wire \line_cache[51][2] ;
 wire \line_cache[51][3] ;
 wire \line_cache[51][4] ;
 wire \line_cache[51][5] ;
 wire \line_cache[51][6] ;
 wire \line_cache[51][7] ;
 wire \line_cache[52][0] ;
 wire \line_cache[52][1] ;
 wire \line_cache[52][2] ;
 wire \line_cache[52][3] ;
 wire \line_cache[52][4] ;
 wire \line_cache[52][5] ;
 wire \line_cache[52][6] ;
 wire \line_cache[52][7] ;
 wire \line_cache[53][0] ;
 wire \line_cache[53][1] ;
 wire \line_cache[53][2] ;
 wire \line_cache[53][3] ;
 wire \line_cache[53][4] ;
 wire \line_cache[53][5] ;
 wire \line_cache[53][6] ;
 wire \line_cache[53][7] ;
 wire \line_cache[54][0] ;
 wire \line_cache[54][1] ;
 wire \line_cache[54][2] ;
 wire \line_cache[54][3] ;
 wire \line_cache[54][4] ;
 wire \line_cache[54][5] ;
 wire \line_cache[54][6] ;
 wire \line_cache[54][7] ;
 wire \line_cache[55][0] ;
 wire \line_cache[55][1] ;
 wire \line_cache[55][2] ;
 wire \line_cache[55][3] ;
 wire \line_cache[55][4] ;
 wire \line_cache[55][5] ;
 wire \line_cache[55][6] ;
 wire \line_cache[55][7] ;
 wire \line_cache[56][0] ;
 wire \line_cache[56][1] ;
 wire \line_cache[56][2] ;
 wire \line_cache[56][3] ;
 wire \line_cache[56][4] ;
 wire \line_cache[56][5] ;
 wire \line_cache[56][6] ;
 wire \line_cache[56][7] ;
 wire \line_cache[57][0] ;
 wire \line_cache[57][1] ;
 wire \line_cache[57][2] ;
 wire \line_cache[57][3] ;
 wire \line_cache[57][4] ;
 wire \line_cache[57][5] ;
 wire \line_cache[57][6] ;
 wire \line_cache[57][7] ;
 wire \line_cache[58][0] ;
 wire \line_cache[58][1] ;
 wire \line_cache[58][2] ;
 wire \line_cache[58][3] ;
 wire \line_cache[58][4] ;
 wire \line_cache[58][5] ;
 wire \line_cache[58][6] ;
 wire \line_cache[58][7] ;
 wire \line_cache[59][0] ;
 wire \line_cache[59][1] ;
 wire \line_cache[59][2] ;
 wire \line_cache[59][3] ;
 wire \line_cache[59][4] ;
 wire \line_cache[59][5] ;
 wire \line_cache[59][6] ;
 wire \line_cache[59][7] ;
 wire \line_cache[5][0] ;
 wire \line_cache[5][1] ;
 wire \line_cache[5][2] ;
 wire \line_cache[5][3] ;
 wire \line_cache[5][4] ;
 wire \line_cache[5][5] ;
 wire \line_cache[5][6] ;
 wire \line_cache[5][7] ;
 wire \line_cache[60][0] ;
 wire \line_cache[60][1] ;
 wire \line_cache[60][2] ;
 wire \line_cache[60][3] ;
 wire \line_cache[60][4] ;
 wire \line_cache[60][5] ;
 wire \line_cache[60][6] ;
 wire \line_cache[60][7] ;
 wire \line_cache[61][0] ;
 wire \line_cache[61][1] ;
 wire \line_cache[61][2] ;
 wire \line_cache[61][3] ;
 wire \line_cache[61][4] ;
 wire \line_cache[61][5] ;
 wire \line_cache[61][6] ;
 wire \line_cache[61][7] ;
 wire \line_cache[62][0] ;
 wire \line_cache[62][1] ;
 wire \line_cache[62][2] ;
 wire \line_cache[62][3] ;
 wire \line_cache[62][4] ;
 wire \line_cache[62][5] ;
 wire \line_cache[62][6] ;
 wire \line_cache[62][7] ;
 wire \line_cache[63][0] ;
 wire \line_cache[63][1] ;
 wire \line_cache[63][2] ;
 wire \line_cache[63][3] ;
 wire \line_cache[63][4] ;
 wire \line_cache[63][5] ;
 wire \line_cache[63][6] ;
 wire \line_cache[63][7] ;
 wire \line_cache[64][0] ;
 wire \line_cache[64][1] ;
 wire \line_cache[64][2] ;
 wire \line_cache[64][3] ;
 wire \line_cache[64][4] ;
 wire \line_cache[64][5] ;
 wire \line_cache[64][6] ;
 wire \line_cache[64][7] ;
 wire \line_cache[65][0] ;
 wire \line_cache[65][1] ;
 wire \line_cache[65][2] ;
 wire \line_cache[65][3] ;
 wire \line_cache[65][4] ;
 wire \line_cache[65][5] ;
 wire \line_cache[65][6] ;
 wire \line_cache[65][7] ;
 wire \line_cache[66][0] ;
 wire \line_cache[66][1] ;
 wire \line_cache[66][2] ;
 wire \line_cache[66][3] ;
 wire \line_cache[66][4] ;
 wire \line_cache[66][5] ;
 wire \line_cache[66][6] ;
 wire \line_cache[66][7] ;
 wire \line_cache[67][0] ;
 wire \line_cache[67][1] ;
 wire \line_cache[67][2] ;
 wire \line_cache[67][3] ;
 wire \line_cache[67][4] ;
 wire \line_cache[67][5] ;
 wire \line_cache[67][6] ;
 wire \line_cache[67][7] ;
 wire \line_cache[68][0] ;
 wire \line_cache[68][1] ;
 wire \line_cache[68][2] ;
 wire \line_cache[68][3] ;
 wire \line_cache[68][4] ;
 wire \line_cache[68][5] ;
 wire \line_cache[68][6] ;
 wire \line_cache[68][7] ;
 wire \line_cache[69][0] ;
 wire \line_cache[69][1] ;
 wire \line_cache[69][2] ;
 wire \line_cache[69][3] ;
 wire \line_cache[69][4] ;
 wire \line_cache[69][5] ;
 wire \line_cache[69][6] ;
 wire \line_cache[69][7] ;
 wire \line_cache[6][0] ;
 wire \line_cache[6][1] ;
 wire \line_cache[6][2] ;
 wire \line_cache[6][3] ;
 wire \line_cache[6][4] ;
 wire \line_cache[6][5] ;
 wire \line_cache[6][6] ;
 wire \line_cache[6][7] ;
 wire \line_cache[70][0] ;
 wire \line_cache[70][1] ;
 wire \line_cache[70][2] ;
 wire \line_cache[70][3] ;
 wire \line_cache[70][4] ;
 wire \line_cache[70][5] ;
 wire \line_cache[70][6] ;
 wire \line_cache[70][7] ;
 wire \line_cache[71][0] ;
 wire \line_cache[71][1] ;
 wire \line_cache[71][2] ;
 wire \line_cache[71][3] ;
 wire \line_cache[71][4] ;
 wire \line_cache[71][5] ;
 wire \line_cache[71][6] ;
 wire \line_cache[71][7] ;
 wire \line_cache[72][0] ;
 wire \line_cache[72][1] ;
 wire \line_cache[72][2] ;
 wire \line_cache[72][3] ;
 wire \line_cache[72][4] ;
 wire \line_cache[72][5] ;
 wire \line_cache[72][6] ;
 wire \line_cache[72][7] ;
 wire \line_cache[73][0] ;
 wire \line_cache[73][1] ;
 wire \line_cache[73][2] ;
 wire \line_cache[73][3] ;
 wire \line_cache[73][4] ;
 wire \line_cache[73][5] ;
 wire \line_cache[73][6] ;
 wire \line_cache[73][7] ;
 wire \line_cache[74][0] ;
 wire \line_cache[74][1] ;
 wire \line_cache[74][2] ;
 wire \line_cache[74][3] ;
 wire \line_cache[74][4] ;
 wire \line_cache[74][5] ;
 wire \line_cache[74][6] ;
 wire \line_cache[74][7] ;
 wire \line_cache[75][0] ;
 wire \line_cache[75][1] ;
 wire \line_cache[75][2] ;
 wire \line_cache[75][3] ;
 wire \line_cache[75][4] ;
 wire \line_cache[75][5] ;
 wire \line_cache[75][6] ;
 wire \line_cache[75][7] ;
 wire \line_cache[76][0] ;
 wire \line_cache[76][1] ;
 wire \line_cache[76][2] ;
 wire \line_cache[76][3] ;
 wire \line_cache[76][4] ;
 wire \line_cache[76][5] ;
 wire \line_cache[76][6] ;
 wire \line_cache[76][7] ;
 wire \line_cache[77][0] ;
 wire \line_cache[77][1] ;
 wire \line_cache[77][2] ;
 wire \line_cache[77][3] ;
 wire \line_cache[77][4] ;
 wire \line_cache[77][5] ;
 wire \line_cache[77][6] ;
 wire \line_cache[77][7] ;
 wire \line_cache[78][0] ;
 wire \line_cache[78][1] ;
 wire \line_cache[78][2] ;
 wire \line_cache[78][3] ;
 wire \line_cache[78][4] ;
 wire \line_cache[78][5] ;
 wire \line_cache[78][6] ;
 wire \line_cache[78][7] ;
 wire \line_cache[79][0] ;
 wire \line_cache[79][1] ;
 wire \line_cache[79][2] ;
 wire \line_cache[79][3] ;
 wire \line_cache[79][4] ;
 wire \line_cache[79][5] ;
 wire \line_cache[79][6] ;
 wire \line_cache[79][7] ;
 wire \line_cache[7][0] ;
 wire \line_cache[7][1] ;
 wire \line_cache[7][2] ;
 wire \line_cache[7][3] ;
 wire \line_cache[7][4] ;
 wire \line_cache[7][5] ;
 wire \line_cache[7][6] ;
 wire \line_cache[7][7] ;
 wire \line_cache[80][0] ;
 wire \line_cache[80][1] ;
 wire \line_cache[80][2] ;
 wire \line_cache[80][3] ;
 wire \line_cache[80][4] ;
 wire \line_cache[80][5] ;
 wire \line_cache[80][6] ;
 wire \line_cache[80][7] ;
 wire \line_cache[81][0] ;
 wire \line_cache[81][1] ;
 wire \line_cache[81][2] ;
 wire \line_cache[81][3] ;
 wire \line_cache[81][4] ;
 wire \line_cache[81][5] ;
 wire \line_cache[81][6] ;
 wire \line_cache[81][7] ;
 wire \line_cache[82][0] ;
 wire \line_cache[82][1] ;
 wire \line_cache[82][2] ;
 wire \line_cache[82][3] ;
 wire \line_cache[82][4] ;
 wire \line_cache[82][5] ;
 wire \line_cache[82][6] ;
 wire \line_cache[82][7] ;
 wire \line_cache[83][0] ;
 wire \line_cache[83][1] ;
 wire \line_cache[83][2] ;
 wire \line_cache[83][3] ;
 wire \line_cache[83][4] ;
 wire \line_cache[83][5] ;
 wire \line_cache[83][6] ;
 wire \line_cache[83][7] ;
 wire \line_cache[84][0] ;
 wire \line_cache[84][1] ;
 wire \line_cache[84][2] ;
 wire \line_cache[84][3] ;
 wire \line_cache[84][4] ;
 wire \line_cache[84][5] ;
 wire \line_cache[84][6] ;
 wire \line_cache[84][7] ;
 wire \line_cache[85][0] ;
 wire \line_cache[85][1] ;
 wire \line_cache[85][2] ;
 wire \line_cache[85][3] ;
 wire \line_cache[85][4] ;
 wire \line_cache[85][5] ;
 wire \line_cache[85][6] ;
 wire \line_cache[85][7] ;
 wire \line_cache[86][0] ;
 wire \line_cache[86][1] ;
 wire \line_cache[86][2] ;
 wire \line_cache[86][3] ;
 wire \line_cache[86][4] ;
 wire \line_cache[86][5] ;
 wire \line_cache[86][6] ;
 wire \line_cache[86][7] ;
 wire \line_cache[87][0] ;
 wire \line_cache[87][1] ;
 wire \line_cache[87][2] ;
 wire \line_cache[87][3] ;
 wire \line_cache[87][4] ;
 wire \line_cache[87][5] ;
 wire \line_cache[87][6] ;
 wire \line_cache[87][7] ;
 wire \line_cache[88][0] ;
 wire \line_cache[88][1] ;
 wire \line_cache[88][2] ;
 wire \line_cache[88][3] ;
 wire \line_cache[88][4] ;
 wire \line_cache[88][5] ;
 wire \line_cache[88][6] ;
 wire \line_cache[88][7] ;
 wire \line_cache[89][0] ;
 wire \line_cache[89][1] ;
 wire \line_cache[89][2] ;
 wire \line_cache[89][3] ;
 wire \line_cache[89][4] ;
 wire \line_cache[89][5] ;
 wire \line_cache[89][6] ;
 wire \line_cache[89][7] ;
 wire \line_cache[8][0] ;
 wire \line_cache[8][1] ;
 wire \line_cache[8][2] ;
 wire \line_cache[8][3] ;
 wire \line_cache[8][4] ;
 wire \line_cache[8][5] ;
 wire \line_cache[8][6] ;
 wire \line_cache[8][7] ;
 wire \line_cache[90][0] ;
 wire \line_cache[90][1] ;
 wire \line_cache[90][2] ;
 wire \line_cache[90][3] ;
 wire \line_cache[90][4] ;
 wire \line_cache[90][5] ;
 wire \line_cache[90][6] ;
 wire \line_cache[90][7] ;
 wire \line_cache[91][0] ;
 wire \line_cache[91][1] ;
 wire \line_cache[91][2] ;
 wire \line_cache[91][3] ;
 wire \line_cache[91][4] ;
 wire \line_cache[91][5] ;
 wire \line_cache[91][6] ;
 wire \line_cache[91][7] ;
 wire \line_cache[92][0] ;
 wire \line_cache[92][1] ;
 wire \line_cache[92][2] ;
 wire \line_cache[92][3] ;
 wire \line_cache[92][4] ;
 wire \line_cache[92][5] ;
 wire \line_cache[92][6] ;
 wire \line_cache[92][7] ;
 wire \line_cache[93][0] ;
 wire \line_cache[93][1] ;
 wire \line_cache[93][2] ;
 wire \line_cache[93][3] ;
 wire \line_cache[93][4] ;
 wire \line_cache[93][5] ;
 wire \line_cache[93][6] ;
 wire \line_cache[93][7] ;
 wire \line_cache[94][0] ;
 wire \line_cache[94][1] ;
 wire \line_cache[94][2] ;
 wire \line_cache[94][3] ;
 wire \line_cache[94][4] ;
 wire \line_cache[94][5] ;
 wire \line_cache[94][6] ;
 wire \line_cache[94][7] ;
 wire \line_cache[95][0] ;
 wire \line_cache[95][1] ;
 wire \line_cache[95][2] ;
 wire \line_cache[95][3] ;
 wire \line_cache[95][4] ;
 wire \line_cache[95][5] ;
 wire \line_cache[95][6] ;
 wire \line_cache[95][7] ;
 wire \line_cache[96][0] ;
 wire \line_cache[96][1] ;
 wire \line_cache[96][2] ;
 wire \line_cache[96][3] ;
 wire \line_cache[96][4] ;
 wire \line_cache[96][5] ;
 wire \line_cache[96][6] ;
 wire \line_cache[96][7] ;
 wire \line_cache[97][0] ;
 wire \line_cache[97][1] ;
 wire \line_cache[97][2] ;
 wire \line_cache[97][3] ;
 wire \line_cache[97][4] ;
 wire \line_cache[97][5] ;
 wire \line_cache[97][6] ;
 wire \line_cache[97][7] ;
 wire \line_cache[98][0] ;
 wire \line_cache[98][1] ;
 wire \line_cache[98][2] ;
 wire \line_cache[98][3] ;
 wire \line_cache[98][4] ;
 wire \line_cache[98][5] ;
 wire \line_cache[98][6] ;
 wire \line_cache[98][7] ;
 wire \line_cache[99][0] ;
 wire \line_cache[99][1] ;
 wire \line_cache[99][2] ;
 wire \line_cache[99][3] ;
 wire \line_cache[99][4] ;
 wire \line_cache[99][5] ;
 wire \line_cache[99][6] ;
 wire \line_cache[99][7] ;
 wire \line_cache[9][0] ;
 wire \line_cache[9][1] ;
 wire \line_cache[9][2] ;
 wire \line_cache[9][3] ;
 wire \line_cache[9][4] ;
 wire \line_cache[9][5] ;
 wire \line_cache[9][6] ;
 wire \line_cache[9][7] ;
 wire \line_cache_idx[2] ;
 wire \line_cache_idx[3] ;
 wire \line_cache_idx[4] ;
 wire \line_cache_idx[5] ;
 wire \line_cache_idx[6] ;
 wire \line_cache_idx[7] ;
 wire \line_cache_idx[8] ;
 wire \line_cache_idx[9] ;
 wire \line_double_counter[0] ;
 wire \line_double_counter[1] ;
 wire \line_double_counter[2] ;
 wire \line_double_counter[3] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net303;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net38;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net39;
 wire net390;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net391;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net392;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net393;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net394;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net395;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net396;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net397;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net398;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net399;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4;
 wire net40;
 wire net400;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \pixel_double_counter[0] ;
 wire \pixel_double_counter[1] ;
 wire \pixel_double_counter[2] ;
 wire \pixel_double_counter[3] ;
 wire \prescaler[0] ;
 wire \prescaler[1] ;
 wire \prescaler[2] ;
 wire \prescaler[3] ;
 wire \prescaler_counter[0] ;
 wire \prescaler_counter[1] ;
 wire \prescaler_counter[2] ;
 wire \prescaler_counter[3] ;
 wire \prescaler_counter[4] ;
 wire \prescaler_counter[5] ;
 wire \prescaler_counter[6] ;
 wire \prescaler_counter[7] ;
 wire \prescaler_counter[8] ;
 wire \res_h_active[0] ;
 wire \res_h_active[1] ;
 wire \res_h_active[2] ;
 wire \res_h_active[3] ;
 wire \res_h_active[4] ;
 wire \res_h_active[5] ;
 wire \res_h_active[6] ;
 wire \res_h_active[7] ;
 wire \res_h_active[8] ;
 wire \res_h_counter[0] ;
 wire \res_h_counter[1] ;
 wire \res_h_counter[2] ;
 wire \res_h_counter[3] ;
 wire \res_h_counter[4] ;
 wire \res_h_counter[5] ;
 wire \res_h_counter[6] ;
 wire \res_h_counter[7] ;
 wire \res_h_counter[8] ;
 wire \res_h_counter[9] ;
 wire \res_v_active[0] ;
 wire \res_v_active[1] ;
 wire \res_v_active[2] ;
 wire \res_v_active[3] ;
 wire \res_v_active[4] ;
 wire \res_v_active[5] ;
 wire \res_v_active[6] ;
 wire \res_v_active[7] ;
 wire \res_v_counter[0] ;
 wire \res_v_counter[1] ;
 wire \res_v_counter[2] ;
 wire \res_v_counter[3] ;
 wire \res_v_counter[4] ;
 wire \res_v_counter[5] ;
 wire \res_v_counter[6] ;
 wire \res_v_counter[7] ;
 wire \res_v_counter[8] ;
 wire \res_v_counter[9] ;
 wire \resolution[0] ;
 wire \resolution[1] ;
 wire \resolution[2] ;
 wire \resolution[3] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_11024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_11551_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_11621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_11621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_11621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_11926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_10408_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_10613_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_10613_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_10148_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_11413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_11413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_11413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_10613_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_10877_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__A (.DIODE(_08848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__C (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A (.DIODE(\res_h_active[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__B (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13257__A (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13257__B (.DIODE(\res_h_active[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__A (.DIODE(\res_h_active[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__B (.DIODE(\res_h_active[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__A (.DIODE(\res_h_active[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__B (.DIODE(\res_h_active[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__A (.DIODE(\res_h_active[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__A (.DIODE(\res_h_active[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__A (.DIODE(\res_h_active[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__B (.DIODE(net3970));
 sky130_fd_sc_hd__diode_2 ANTENNA__13274__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__A (.DIODE(\res_h_active[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13278__B (.DIODE(\res_h_active[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__A1 (.DIODE(\res_h_active[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13282__A (.DIODE(\res_h_active[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__B (.DIODE(\res_h_active[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13287__B (.DIODE(\res_h_active[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__B (.DIODE(\res_h_active[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13301__B (.DIODE(\res_h_active[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__A1 (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13313__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13315__A (.DIODE(_08848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__B1 (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__A (.DIODE(\res_h_active[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A (.DIODE(\res_h_active[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A (.DIODE(net3966));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__B (.DIODE(net3966));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__A (.DIODE(net3971));
 sky130_fd_sc_hd__diode_2 ANTENNA__13334__B (.DIODE(net3971));
 sky130_fd_sc_hd__diode_2 ANTENNA__13340__B (.DIODE(\res_h_active[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13342__A (.DIODE(\res_h_active[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13342__B (.DIODE(\res_h_active[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__B1 (.DIODE(\res_h_active[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__B (.DIODE(\res_h_active[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13357__B1 (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__A1 (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__A (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__13369__A (.DIODE(_09107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13371__A (.DIODE(_09105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13371__B (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__B (.DIODE(_09111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13373__A (.DIODE(_09105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13375__A (.DIODE(_08848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__B (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__A1 (.DIODE(_09112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__B (.DIODE(_08848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__C (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__B (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__B1 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__B2 (.DIODE(_08848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__B (.DIODE(_09112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__A (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__C (.DIODE(_09128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A2 (.DIODE(_09105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__A1 (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13760__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A (.DIODE(_08848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__B (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__A (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__A (.DIODE(_09498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13769__C (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__C (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__B (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13782__A (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13788__B (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13793__B (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__A (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__B (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__A (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__A (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13806__A (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13808__B (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__B (.DIODE(_09536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13812__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13815__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13817__A (.DIODE(_09542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__B (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__A (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__A (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__A (.DIODE(_09549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13825__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13828__A (.DIODE(_09553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13833__A (.DIODE(_09558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13834__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13834__B (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13838__A (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13839__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13839__B (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13843__A (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13843__B (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13844__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13844__B (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__C (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13848__C (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13852__A (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13852__B (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13854__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13854__B (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13854__C (.DIODE(_09579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13856__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13856__B (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__A (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__B (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__A1 (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__A2 (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__B (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__A (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__B (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__A (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__B (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13870__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__D (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__A (.DIODE(_09600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__B (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13880__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13880__B (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13882__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13882__B (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13884__B (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13885__A (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13886__B1 (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__A2 (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__A1 (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__A2 (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__B1 (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13890__A (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__A (.DIODE(_09542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__A (.DIODE(_09617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__A (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A (.DIODE(_09617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__B (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__C (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__A (.DIODE(_09624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A (.DIODE(_09626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13906__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13906__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__B (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13909__C (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__B (.DIODE(_09637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__C (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__A (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__B (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__A (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__B (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13917__A (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__B (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__C (.DIODE(_09643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__B (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__C (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__A (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A (.DIODE(_09650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__B (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__C (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__B (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__C (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__B (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__C (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13936__A (.DIODE(_09579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__B (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__C (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__A (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__B (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__C (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13938__D (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__A (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__B (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13939__C (.DIODE(_09653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__A (.DIODE(_09536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13941__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13943__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13943__B (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__A (.DIODE(_09553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13946__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__B (.DIODE(_09673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13950__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13950__B (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13950__C (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__B (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__C (.DIODE(_09558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__B (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13952__C (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13953__A (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13953__B (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__A (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__B (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__B (.DIODE(_09681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13956__C (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__B (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__C (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13960__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__A (.DIODE(_09687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__A (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13966__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__A (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__B (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__C (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__D (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__B (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__C (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__B (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13972__C (.DIODE(_09643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__A (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__A (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__A1 (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13978__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13978__B (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13978__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__B (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__C (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__B (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__C (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__B (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__C (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__A (.DIODE(_09549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__A (.DIODE(_09714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__C (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__B (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__B (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__B (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__C (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__A (.DIODE(_09714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__B (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__B (.DIODE(_09637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__B (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__C (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__A1 (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__B1 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__C1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__D1 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14009__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14011__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__B (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__C (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__B (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__C (.DIODE(_09643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__A (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14019__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14021__A (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14021__B (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A (.DIODE(_09549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__C (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__A (.DIODE(_09751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A (.DIODE(_09542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__C (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14028__A (.DIODE(_09753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__A (.DIODE(_09553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__C (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__A (.DIODE(_09755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__A (.DIODE(_09536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__C (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__A (.DIODE(_09757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__A1 (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__A3 (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__A4 (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__B1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14036__A (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14036__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__A (.DIODE(_09542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14038__A (.DIODE(_09763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__A (.DIODE(_09549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14040__B (.DIODE(_09536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__B (.DIODE(_09553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14042__A (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__A1 (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__A2 (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__A3 (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__A4 (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__B1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__C (.DIODE(_09770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__A (.DIODE(_09714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__B (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14046__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14048__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14048__B (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14048__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14050__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14051__A (.DIODE(_09776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__B (.DIODE(_09637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__C (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__B (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__C (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__D (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__A (.DIODE(_09714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__B (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__C (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__B (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__B (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__C (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__B (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__C (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__A (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__B (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__C (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__D (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14065__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__A (.DIODE(_09791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14067__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__A (.DIODE(_09793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__A (.DIODE(_09795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14071__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__A (.DIODE(_09797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__A (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__B (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__C (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14073__D (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__B (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__C (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14076__A (.DIODE(_09715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14076__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14076__C (.DIODE(_09643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14078__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14078__B (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14079__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__A (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__C (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__B (.DIODE(_09681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__C (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__C (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__A (.DIODE(_09812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__A (.DIODE(_09687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__A (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__B (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__C (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14090__D (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__B (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__C (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14092__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14092__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14092__C (.DIODE(_09643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14094__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14096__A (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__B (.DIODE(_09673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__C (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__C (.DIODE(_09568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__C (.DIODE(_09558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__B (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__C (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14103__D (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14104__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14104__B (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14104__C (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14105__A (.DIODE(_09671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14105__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14105__C (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__B (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__C (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__A (.DIODE(_09672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__C (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14111__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14115__A3 (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14115__B1 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__B (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__C (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14123__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14123__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14125__C (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14126__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14126__B (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__B (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14130__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14130__C (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__B (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__C (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__D (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__A (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14139__A (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__A (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14143__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14145__A (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14146__A (.DIODE(_09871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14146__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14148__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14148__B (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14148__C (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14148__D (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14149__A (.DIODE(_09841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__B (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14150__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14152__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14152__B (.DIODE(_09558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14152__C (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14153__A (.DIODE(_09624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14153__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__A (.DIODE(_09626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__A (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__B (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__B (.DIODE(_09637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14159__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14159__B (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14159__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14161__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14161__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14161__C (.DIODE(_09681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14163__A1 (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14163__A2 (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14164__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14164__B (.DIODE(_09656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14164__C (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14165__A (.DIODE(_09617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14165__B (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14168__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14170__A (.DIODE(_09621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14170__B (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14170__C (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14171__A (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14171__B (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14171__C (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14171__D (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14173__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14175__A (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14178__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14180__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__A (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__B (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__C (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14186__A (.DIODE(_09771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14187__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14187__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14194__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14194__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14195__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14197__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14198__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14200__A (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14203__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14207__B1 (.DIODE(\line_cache[287][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14209__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14221__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14221__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14224__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14224__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14227__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14227__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14228__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14229__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14229__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14237__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14239__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14239__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14245__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14245__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14248__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14248__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14250__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14250__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14251__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14251__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14252__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14252__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14253__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14253__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14255__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14257__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14257__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14260__B (.DIODE(_09957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14266__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14266__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14268__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14268__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14271__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14271__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14272__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14272__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14272__C (.DIODE(_09662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14273__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14273__B (.DIODE(_09659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14273__C (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14275__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14275__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__B (.DIODE(_09577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__C (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14278__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__B (.DIODE(_09634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14280__C (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14283__A (.DIODE(_09668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14283__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14283__C (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14291__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14293__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14293__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14294__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14302__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14302__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14304__B (.DIODE(_10029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__B (.DIODE(_09607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14306__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14311__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14311__B (.DIODE(_09605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__A (.DIODE(_09646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__B (.DIODE(_09530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__A (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14316__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__A (.DIODE(_10044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14320__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14320__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14321__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14321__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14322__A (.DIODE(_09563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14324__A (.DIODE(_09681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14324__B (.DIODE(_08995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14325__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14325__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14328__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14329__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14330__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14330__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14331__A (.DIODE(_09541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14331__B (.DIODE(_09579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14332__A (.DIODE(_10057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14333__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14333__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14334__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14334__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14335__A (.DIODE(_08993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14336__A (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__A (.DIODE(_09537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__A (.DIODE(_09650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14341__A (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14342__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14343__A (.DIODE(_09673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14344__A (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14346__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__A (.DIODE(_09558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__B (.DIODE(_09778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__A (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14350__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14350__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14353__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14353__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14359__B (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14361__A (.DIODE(_09871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14361__B (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14364__C1 (.DIODE(_10089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__A1 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14366__A1 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14366__B2 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14367__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14367__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14368__A1 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14368__B2 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14372__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14375__A (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14376__A (.DIODE(_10044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14377__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14378__A (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14380__A (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14381__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__A (.DIODE(_09600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14385__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14386__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14387__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14392__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14392__B (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14394__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14394__B (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14398__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14398__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__A (.DIODE(_09550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14405__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14405__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__B (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14407__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14407__B (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14410__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14410__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14411__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14411__B (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__B (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__B (.DIODE(_09616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14414__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14416__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14416__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14417__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14417__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14418__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14418__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14419__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14419__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14422__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14422__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14426__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14426__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14428__A (.DIODE(_09543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14428__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14433__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14433__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14434__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14438__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14438__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14442__A (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14442__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14442__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14443__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14443__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14444__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14444__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__B (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14449__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14449__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14450__A (.DIODE(_10057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14451__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14451__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14454__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14454__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14455__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14455__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__B (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__B (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14461__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14461__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14462__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14462__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__B (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14464__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14464__B (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14467__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14467__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14470__A (.DIODE(_09555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14470__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14473__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14473__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14474__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14474__B (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14480__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14480__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14485__A (.DIODE(_09554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14485__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__A (.DIODE(_10192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14489__A (.DIODE(_10186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14490__C (.DIODE(_10158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14490__D (.DIODE(_10215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14491__A (.DIODE(_09753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14491__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14491__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__A (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__A (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__A (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14497__A (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14498__A (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__A (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14500__A (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__A (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14504__A (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14505__A (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14506__A (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__A (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14510__A (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14511__A (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14512__A (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__A (.DIODE(_09751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__A (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__A (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__A (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14520__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14522__A (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14522__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14523__A (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14523__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__A (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14525__A (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14525__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14528__A (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14528__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14529__A (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14529__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__A (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__A (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14531__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__A (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__A (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__A (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__B (.DIODE(_09752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14541__A (.DIODE(_09551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14541__B (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__A (.DIODE(_10267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14543__A (.DIODE(_10268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14543__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__A (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__A (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14549__A (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14549__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__A (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__A (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__A (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14552__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14555__B (.DIODE(_10280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__A (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__A (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14559__A (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14559__B (.DIODE(_09756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__A (.DIODE(_09755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__C (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__A3 (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14567__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14570__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14570__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14571__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14571__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__B (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__B (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14576__A (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14577__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14577__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14578__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14578__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__B (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14583__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14583__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14585__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14585__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14586__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14586__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14589__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14589__B (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14590__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14591__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14591__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__A (.DIODE(_09768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14595__A (.DIODE(_10301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__A (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__A (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14598__A (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14602__A (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14602__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14603__A (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14603__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__A (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__C (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__A (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__B (.DIODE(_10268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14609__A (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14609__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14610__A (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14610__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14611__A (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14611__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14613__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__A (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__A (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__A (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__A (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14625__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14625__B (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14626__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14626__B (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14629__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14631__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__A (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14638__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14638__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14639__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14639__B (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14640__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14640__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14642__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14643__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14643__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14644__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14644__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14645__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14645__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__A (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__A (.DIODE(_10354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__B (.DIODE(_10048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14651__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14651__B (.DIODE(_10073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__B (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14653__B (.DIODE(_09569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__A (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__B (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__C (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14657__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14657__B (.DIODE(_10115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__B (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14659__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14659__B (.DIODE(_10032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__B (.DIODE(_10062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14663__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14663__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__A (.DIODE(_09763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__B (.DIODE(_10050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14665__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14665__B (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__B (.DIODE(_10119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14669__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14669__B (.DIODE(_10055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14670__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14670__B (.DIODE(_09578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14671__A (.DIODE(_09764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14671__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__A (.DIODE(_10381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A (.DIODE(_10295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__C (.DIODE(_10401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14677__B (.DIODE(_10216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14677__C (.DIODE(_10402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14678__A2 (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14679__A (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14680__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14681__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14681__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14686__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14699__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14704__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14708__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14710__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14710__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14711__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14711__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14713__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14715__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14715__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14717__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14718__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14738__A (.DIODE(_10418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14738__C (.DIODE(_10462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14739__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14740__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14740__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14741__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14741__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14749__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14749__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__C1 (.DIODE(_10479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__A1 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__B2 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14757__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14758__A1 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14758__B2 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14759__A2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14759__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14769__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14769__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14770__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14770__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14780__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14780__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14782__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14782__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14783__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14789__B (.DIODE(_10513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14790__A (.DIODE(_10487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14791__A (.DIODE(_10463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14794__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14794__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14795__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14795__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14796__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14797__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14798__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14803__B1 (.DIODE(\line_cache[287][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14807__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14808__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14810__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14810__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14820__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14820__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14823__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14823__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14825__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14829__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14831__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14831__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14832__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14833__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14835__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14835__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14839__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14839__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14842__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14842__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14843__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14844__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14844__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14845__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14845__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14846__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14846__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14847__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14847__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14848__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14849__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14854__B (.DIODE(_10552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14856__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14859__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14860__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14860__B (.DIODE(_09751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14871__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14872__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14873__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14874__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14877__A_N (.DIODE(_10593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14889__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__A (.DIODE(_09545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__B (.DIODE(_09767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__C (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14897__A (.DIODE(_10621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14900__B (.DIODE(_10618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14901__A (.DIODE(_09596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14901__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14904__A (.DIODE(_10069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14904__B (.DIODE(_09760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14908__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14912__B (.DIODE(_10636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14916__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__14920__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14927__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14933__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14935__C (.DIODE(_10650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14937__A (.DIODE(_10613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14937__C (.DIODE(_10661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__C (.DIODE(_10662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14939__B1_N (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__A (.DIODE(_10664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14945__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14945__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14946__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14946__B (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14948__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14948__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14952__A1 (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14952__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14957__A (.DIODE(_10668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14958__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14958__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14959__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14959__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14960__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14960__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14961__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14964__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14965__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14965__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14967__B (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14968__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14969__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14970__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14976__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14977__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14981__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14981__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14984__C1 (.DIODE(_10707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14985__A1 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14985__B2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14986__A1 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14986__B2 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14987__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14987__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14988__A1 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14988__B2 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14992__A (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14993__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14994__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14997__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14997__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14998__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15000__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15009__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15019__B (.DIODE(_10742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15026__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15026__B (.DIODE(_10045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__A (.DIODE(_09766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__B (.DIODE(_10058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15038__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15043__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15047__A (.DIODE(_10756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15048__D (.DIODE(_10771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15051__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15051__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15052__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15052__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15053__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15054__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15055__A1 (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__B1 (.DIODE(\line_cache[287][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15062__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15064__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15065__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15067__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15067__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15068__C_N (.DIODE(_10791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15081__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15085__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15086__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15088__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15088__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15089__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15092__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15092__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15094__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15094__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15099__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15099__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15100__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15100__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15101__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15101__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15102__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15102__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15103__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15104__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15106__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15106__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15108__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15108__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15109__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15109__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__B (.DIODE(_10808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15119__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15121__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15122__B (.DIODE(_10841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15127__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15133__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15135__C (.DIODE(_10850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15146__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15150__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15160__A (.DIODE(_09755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15160__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15162__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15165__A_N (.DIODE(_10880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15176__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15176__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15179__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15179__C (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15183__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15188__B (.DIODE(_10890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15189__A (.DIODE(_10772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15189__C (.DIODE(_10912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15190__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15191__B1 (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15196__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15196__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15197__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15197__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15198__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15198__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15200__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15200__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15216__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15221__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15221__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15222__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15222__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15223__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15225__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15225__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15227__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15237__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15248__A (.DIODE(_10928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15249__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15250__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15250__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15251__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15251__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15262__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15262__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15265__C1 (.DIODE(_10987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15266__A1 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15266__B2 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15267__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15267__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15268__A1 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15268__B2 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15269__A2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15269__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15277__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15277__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15278__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15278__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15279__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15279__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15282__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15282__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15284__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15284__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15290__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15290__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15292__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15292__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15293__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15296__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15297__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15297__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__B (.DIODE(_11021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__A (.DIODE(_10995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15301__A (.DIODE(_10971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15304__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15304__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15305__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15305__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15306__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15307__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15313__B1 (.DIODE(\line_cache[287][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15318__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15330__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15330__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15333__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15333__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15334__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15335__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15335__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15338__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15339__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15342__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15345__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15345__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15347__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15347__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15349__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15349__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15352__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15352__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15353__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15353__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15354__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15354__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15355__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15355__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15356__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15356__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15358__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15359__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15361__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15361__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15364__B (.DIODE(_11060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15365__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15366__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15369__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__B (.DIODE(_09751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15379__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15380__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15381__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15382__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15400__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15404__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15410__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15411__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15412__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15416__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15418__C (.DIODE(_11132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15420__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15430__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15430__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15433__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15433__B (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15442__A (.DIODE(_11119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15442__B (.DIODE(_11142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15443__C (.DIODE(_11165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15444__B1_N (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15445__A (.DIODE(_11167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15446__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15447__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15447__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15448__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15448__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15449__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15449__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15463__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15468__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15471__A (.DIODE(_11181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15472__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15473__A (.DIODE(_10044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15473__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15474__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15474__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15475__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15477__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15477__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15478__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15479__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15480__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15489__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15500__A (.DIODE(_11179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15501__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15502__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15502__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15503__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15503__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15511__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15511__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15517__C1 (.DIODE(_11238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15518__A1 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15518__B2 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15519__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15519__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__A1 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__B2 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__A2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15530__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15530__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15532__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15532__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15534__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15534__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15536__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15536__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15542__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15542__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15543__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15543__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15544__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15544__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15545__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15548__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__B (.DIODE(_11272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15556__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15556__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15557__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15557__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15558__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15559__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15560__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15565__B1 (.DIODE(\line_cache[287][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15567__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15569__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15570__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15582__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15582__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15585__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15585__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15586__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15587__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15587__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15590__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15591__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15594__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15595__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15606__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15606__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15607__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15607__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15609__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15609__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15613__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15613__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15616__B (.DIODE(_11311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15620__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15630__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15631__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15636__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15638__C (.DIODE(_11351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15640__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15650__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15650__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15658__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15660__B (.DIODE(_11381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15662__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15665__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15669__C (.DIODE(_11388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15674__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15676__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15677__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15680__A_N (.DIODE(_11393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15691__A (.DIODE(_11391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15692__A (.DIODE(_11361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15692__C (.DIODE(_11413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15693__A (.DIODE(_11275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15693__B (.DIODE(_11338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15693__C (.DIODE(_11414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__B1_N (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__A (.DIODE(_11416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15696__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15697__A (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15697__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15700__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15700__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15701__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15701__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15715__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15720__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15724__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15725__A (.DIODE(_10044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15726__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15726__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15727__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15729__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15729__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15730__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15731__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15732__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15741__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15752__A (.DIODE(_11430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15752__C (.DIODE(_11472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15753__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15754__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15754__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15755__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15755__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15761__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15761__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15762__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15762__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15763__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15763__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__C (.DIODE(_11481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15766__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15766__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15770__A1 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15770__B2 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15771__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15771__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15772__A1 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15772__B2 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15773__A2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15773__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15781__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15781__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15782__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15782__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15784__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15784__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15786__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15786__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15795__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15795__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15796__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15796__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15797__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15800__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15801__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15801__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15803__B (.DIODE(_11523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15805__B (.DIODE(_11525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15808__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15808__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15809__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15809__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15810__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15811__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15812__A1 (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15817__B1 (.DIODE(\line_cache[287][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15819__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15821__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15822__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15824__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15824__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15831__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15831__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15834__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15834__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15837__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15837__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15838__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15842__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15843__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15845__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15845__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15846__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15847__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15849__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15849__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15851__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15851__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15853__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15853__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15856__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15856__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15857__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15857__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15859__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15859__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15861__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15861__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15862__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15863__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15868__B (.DIODE(_11562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15873__A (.DIODE(_09753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15873__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15873__D (.DIODE(_09683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15883__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15884__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15885__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15886__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__A_N (.DIODE(_11601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15891__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15894__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15904__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__15908__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15909__A (.DIODE(_11623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15914__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15915__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15920__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15922__C (.DIODE(_11634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15924__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15939__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__B (.DIODE(_11663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15944__A (.DIODE(_11621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15945__B (.DIODE(_11589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15945__C (.DIODE(_11665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15946__B1_N (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15947__A (.DIODE(_11667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15948__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15949__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15949__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15951__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15951__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15965__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15970__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15975__A (.DIODE(_10044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15977__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15979__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15979__C (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15980__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15981__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15982__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15991__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16002__A (.DIODE(_11679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16003__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16004__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16004__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16005__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16005__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16011__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16011__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16013__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16013__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16016__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16016__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16020__A1 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16020__B2 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16021__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16021__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16022__A1 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16022__B2 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16023__A2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16023__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16026__A (.DIODE(_11735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16032__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16032__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16033__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16033__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16046__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16046__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16047__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16050__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16051__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16051__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16053__B (.DIODE(_11772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16055__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16058__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16058__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16059__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16059__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16060__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16061__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16062__A1 (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16067__B1 (.DIODE(\line_cache[287][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16069__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16071__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16072__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16081__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16081__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16087__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16087__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16088__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16089__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16089__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16092__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16093__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16095__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16095__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16096__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16097__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16099__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16099__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16101__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16101__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16103__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16103__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16106__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16106__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16107__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16107__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16108__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16108__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16109__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16109__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16110__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16110__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16111__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16111__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16112__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16113__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16115__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16115__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16116__D (.DIODE(_11835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16118__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16119__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16120__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16123__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16124__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16124__B (.DIODE(_09751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16133__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16134__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16135__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16136__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16153__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16157__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16163__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16164__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16165__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16169__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16171__C (.DIODE(_11882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16173__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16173__B (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16175__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16176__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16176__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16179__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16179__C (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__A (.DIODE(_11869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__B (.DIODE(_11892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16196__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16196__C (.DIODE(_11915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16197__B1_N (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16198__A (.DIODE(_11917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16199__A (.DIODE(_09912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16200__A (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16200__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16201__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16201__C (.DIODE(_10167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16202__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16202__C (.DIODE(_10161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16216__A_N (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16221__A_N (.DIODE(_09597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16225__A (.DIODE(_09595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16226__A (.DIODE(_10044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16227__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16227__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16228__A (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16230__A (.DIODE(_09544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16230__C (.DIODE(_09600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16231__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16232__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16232__C (.DIODE(_10434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16233__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16242__B1 (.DIODE(_10139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16252__B (.DIODE(_11970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16253__A (.DIODE(_11929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16253__C (.DIODE(_11971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16254__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16255__A (.DIODE(_10038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16255__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16256__A (.DIODE(_10041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16256__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16262__A (.DIODE(_10067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16262__C (.DIODE(_10075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16263__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16263__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16264__A (.DIODE(_10074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16264__C (.DIODE(_09540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16267__A1 (.DIODE(_09623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16267__B1 (.DIODE(_09620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16270__C1 (.DIODE(_11988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16271__A1 (.DIODE(_09658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16271__B2 (.DIODE(_09661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16272__A1 (.DIODE(_09645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16272__B2 (.DIODE(_09648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16273__A1 (.DIODE(_09639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16273__B2 (.DIODE(_09636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16274__A2 (.DIODE(_09663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16274__B2 (.DIODE(_09655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__B (.DIODE(_09546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16283__A (.DIODE(_09848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16283__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16284__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16284__B (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16285__A (.DIODE(_09840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16285__B (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16287__A (.DIODE(_09858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16287__B (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16289__A1 (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16289__A3 (.DIODE(_09862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16294__A (.DIODE(_12000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16295__A1 (.DIODE(_09682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16295__B2 (.DIODE(_09685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16296__A2 (.DIODE(_09689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16296__B2 (.DIODE(_09693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16297__A1 (.DIODE(_09728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16297__B2 (.DIODE(_09726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16298__A2 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16301__A1 (.DIODE(_10025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16302__A2 (.DIODE(_10023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16302__B2 (.DIODE(_10024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16304__B (.DIODE(_12022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16306__B (.DIODE(_12024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16309__A (.DIODE(_09917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16309__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16310__A (.DIODE(_09919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16310__B (.DIODE(_09532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16311__A2 (.DIODE(_09867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16312__B (.DIODE(_09531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16313__A1 (.DIODE(_09547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16318__B1 (.DIODE(\line_cache[287][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16320__B2 (.DIODE(_09804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16322__A (.DIODE(_09787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16323__A (.DIODE(_09789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__A1 (.DIODE(_09785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__B2 (.DIODE(_09801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16332__A1 (.DIODE(_09675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16332__B2 (.DIODE(_09676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16335__A1 (.DIODE(_09677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16335__B2 (.DIODE(_09678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16338__A1 (.DIODE(_09809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16338__B2 (.DIODE(_09811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16339__B2 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16340__A1 (.DIODE(_09813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16340__B2 (.DIODE(_09815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16343__A (.DIODE(_09864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16344__A (.DIODE(_09860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16346__A1 (.DIODE(_09870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16346__B2 (.DIODE(_09873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16347__A (.DIODE(_09853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16348__A (.DIODE(_09857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16350__A1 (.DIODE(_09855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16350__B1 (.DIODE(_09847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16352__A (.DIODE(_09631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16352__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16354__A1 (.DIODE(_09877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16354__B2 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16357__A1 (.DIODE(_09796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16357__B2 (.DIODE(_09798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__A2 (.DIODE(_09777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__B2 (.DIODE(_09794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16359__A1 (.DIODE(_09890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16359__B2 (.DIODE(_09896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__A2 (.DIODE(_09892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__B2 (.DIODE(_09895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16361__A1 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16361__B2 (.DIODE(_09900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16362__A2 (.DIODE(_09792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16362__B2 (.DIODE(_09905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16363__A (.DIODE(_09773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16364__A (.DIODE(_09775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16366__A1 (.DIODE(_09783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16366__B2 (.DIODE(_09780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__C_N (.DIODE(_12086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16370__A1 (.DIODE(_10244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16371__A2 (.DIODE(_10242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16374__B2 (.DIODE(_10257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16375__A (.DIODE(_10104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16375__B (.DIODE(_09751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16384__B (.DIODE(_10102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16385__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16386__A3 (.DIODE(_10106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16387__A3 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16405__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__A2 (.DIODE(_10394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16410__A (.DIODE(_12122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__A (.DIODE(_10035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16416__A (.DIODE(_10176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16417__A (.DIODE(_10054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16421__A2 (.DIODE(_10363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16423__C (.DIODE(_12133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16425__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16425__B (.DIODE(_10031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16427__A2 (.DIODE(_10334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__A (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__B (.DIODE(_10098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16431__A (.DIODE(_10071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16431__C (.DIODE(_09758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16445__A (.DIODE(_12157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__A (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__B (.DIODE(_12088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__C (.DIODE(_12166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__B1_N (.DIODE(_08979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16450__A (.DIODE(_12168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16452__A (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16456__B (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16458__A (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16458__B (.DIODE(_12175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16460__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16462__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16463__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16465__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__16466__A (.DIODE(_12183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__A (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16468__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16470__B (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__16472__A (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16473__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16473__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16475__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16478__A (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__16480__A (.DIODE(_12196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__A (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16482__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16484__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16487__A (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16488__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__A (.DIODE(_12204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16490__A (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16491__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16492__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16492__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16493__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16496__A (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16497__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__16498__A (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__A (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16501__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16501__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16502__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16505__A (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16506__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__16507__A (.DIODE(_12220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__A (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16509__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16511__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16514__A (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__16516__A (.DIODE(_12228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16517__A (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16518__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16520__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16523__A (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16524__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__16525__A (.DIODE(_12236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16526__A (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16528__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16528__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16532__A (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16533__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__16534__A (.DIODE(_12244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16535__A (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16536__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16537__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16537__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16538__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16540__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__16540__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__16542__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__16544__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__16547__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__16547__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__16548__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__16549__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__16550__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__16550__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__16552__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__16553__B (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16557__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__16557__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__16558__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__16561__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__16563__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__16563__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16566__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16566__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__16567__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16572__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__16572__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__16575__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__16575__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__16576__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__16579__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__16579__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__16582__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__16587__A (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16588__A (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__B (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__C (.DIODE(_09105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16590__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__A1 (.DIODE(_12292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__A2 (.DIODE(_12293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__B1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16594__A2 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16594__B1 (.DIODE(_09112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16595__B (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16595__C (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16596__A (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16597__A1 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16598__A (.DIODE(_09111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16600__A2 (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__A (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16603__C (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16604__A2 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16604__B1 (.DIODE(_09112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__B (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16608__A (.DIODE(_09111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16610__A2 (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__B (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16613__A (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16614__A1 (.DIODE(_09112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16614__B2 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16616__A1 (.DIODE(_12311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16616__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16616__B1 (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16618__A (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16618__B (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__A (.DIODE(_09111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16623__A (.DIODE(_09111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16633__A (.DIODE(_09107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16635__A (.DIODE(_12326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16635__B (.DIODE(_12328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16637__B (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16640__A (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16641__A2 (.DIODE(_12332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16645__A (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16646__A1 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16646__A2 (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16647__B (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16649__B (.DIODE(_09107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16650__A (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16654__B1 (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16656__A (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16657__B1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__A1 (.DIODE(_12326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__A2 (.DIODE(_12328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__A1 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__B1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16661__A1 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16663__B (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16664__B (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16671__B1 (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16675__B1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16678__A (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16683__B1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16686__A (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16691__B1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16694__A (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16695__B1 (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16698__B1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16701__A (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16705__B1 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16705__C1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16706__B (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16707__A1 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16708__B1 (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16717__A2 (.DIODE(_12332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16717__B2 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16719__B (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16720__A1 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16721__B (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16728__A2 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16729__A2 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16730__A3 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16730__B1 (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16736__A2 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16737__A2 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16738__C (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16739__A (.DIODE(_12342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__A1 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__C1 (.DIODE(_12341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16748__B (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16749__A3 (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16749__A4 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16753__A2 (.DIODE(_12332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16753__B2 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16759__B (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16760__A3 (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16760__A4 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16764__A2 (.DIODE(_12332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16764__B2 (.DIODE(_12337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16769__B (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16770__A3 (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16770__A4 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16774__B (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16775__A2 (.DIODE(_09106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16775__A4 (.DIODE(_12333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16776__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16778__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16780__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16782__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16784__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__16784__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16786__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__16786__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16790__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__16790__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16792__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16794__S (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16796__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16799__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__16799__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16801__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16801__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16807__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__16807__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16809__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__16809__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16811__A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__16811__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16823__A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__16823__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16827__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__16827__S (.DIODE(_12450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16829__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16830__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__16830__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16832__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__16832__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16834__A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__16834__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16836__A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__16836__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16838__A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__16838__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16840__A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__16840__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16842__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__16842__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16844__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__16844__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16846__A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__16846__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16848__A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__16848__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16852__A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__16852__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16854__A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__16854__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16856__A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__16856__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16858__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__16858__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16860__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__16860__S (.DIODE(_12467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16862__A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16862__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16864__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__16864__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16866__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__16866__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16870__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__16870__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16872__A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__16872__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16874__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__16874__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16876__A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__16876__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16884__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__16884__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16886__A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__16886__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16888__A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__16888__S (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16890__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__16890__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__16894__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__16894__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16895__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__16898__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16898__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__16899__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__16902__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__16902__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__16903__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16906__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__16906__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__16907__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__16910__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__16910__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__16911__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__16914__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__16914__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__16915__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__16916__A1 (.DIODE(net3970));
 sky130_fd_sc_hd__diode_2 ANTENNA__16918__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__16918__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__16919__A1 (.DIODE(net3966));
 sky130_fd_sc_hd__diode_2 ANTENNA__16921__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__16922__A1 (.DIODE(net3971));
 sky130_fd_sc_hd__diode_2 ANTENNA__17081__B (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17082__A (.DIODE(_09498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17089__A2 (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17089__B2 (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17091__A2 (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17091__B2 (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17095__A2 (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17095__B2 (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17099__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17099__B2 (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17103__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17103__B2 (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17107__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17107__B2 (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17112__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17116__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17118__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17119__A (.DIODE(\base_v_bporch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17121__B (.DIODE(\base_v_bporch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17130__B (.DIODE(\base_v_bporch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17131__B1 (.DIODE(\base_v_bporch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17237__B (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__17243__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__17244__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__17245__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17247__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17247__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17248__B (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17249__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17252__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17254__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17255__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17257__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__17257__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__17258__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__17258__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__17260__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__17263__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17264__B (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17267__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17267__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17268__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17273__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17274__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17275__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__17277__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__17277__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__17278__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__17278__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__17287__B (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17290__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17290__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17291__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17296__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17297__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__B (.DIODE(_12885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17301__A (.DIODE(_12885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17306__B1 (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17308__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17308__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17309__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17313__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17315__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17317__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__17318__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__17319__B (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17321__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17321__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17322__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17326__A (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17328__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17330__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17334__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17338__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17340__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17341__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__17342__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__17344__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17346__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17346__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17347__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17351__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17353__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17354__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__17356__A (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17357__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__17359__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17359__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17360__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17364__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17365__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17367__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__17367__B1 (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17370__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17370__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17371__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17373__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17375__A (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17376__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17378__B (.DIODE(_12686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17378__C (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17379__A (.DIODE(_12837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17382__A (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17382__B (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17384__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17385__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__17393__A (.DIODE(_12971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17396__C1 (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17401__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17402__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17402__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17406__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17406__C (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17407__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17407__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17410__B (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17411__B (.DIODE(_09601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17417__A (.DIODE(_10109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17417__B (.DIODE(_09553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17418__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17419__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17419__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17422__A (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17423__B (.DIODE(_09013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17424__B (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17425__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17425__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17427__A2 (.DIODE(_12971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17429__B (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17430__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17430__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17432__A2 (.DIODE(_12971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17433__B (.DIODE(_09533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17434__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17435__B (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17436__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17436__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17437__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17438__A2 (.DIODE(_12971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17440__B1 (.DIODE(_09127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17441__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17443__A2 (.DIODE(_12971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17445__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17445__B (.DIODE(_12825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17490__B1 (.DIODE(_09516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17491__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17512__A (.DIODE(_09498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17518__A_N (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17523__A (.DIODE(_13085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17524__A2 (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17531__A (.DIODE(_13085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17532__A2 (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17538__A (.DIODE(_09498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17546__A (.DIODE(_13085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17547__A2 (.DIODE(_12682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17553__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17559__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17566__A2 (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17572__A (.DIODE(_13085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17573__A (.DIODE(_09498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17576__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17577__B (.DIODE(_09497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17583__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17589__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17592__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17594__A (.DIODE(_12960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__B (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17599__B (.DIODE(_09052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17613__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17613__B (.DIODE(_12183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17615__A (.DIODE(_02809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17620__A (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17622__A (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17623__A (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17624__A1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17624__A2 (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17624__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17625__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17625__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17627__A (.DIODE(_09126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17627__B (.DIODE(_12196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17629__A (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17630__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17630__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17632__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17632__B (.DIODE(_12204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17634__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17635__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17635__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17637__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17637__B (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17639__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17640__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17640__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__B (.DIODE(_12220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17644__A (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17645__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17645__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17647__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17647__B (.DIODE(_12228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17649__A (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17650__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17650__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17652__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17652__B (.DIODE(_12236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17654__A (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17655__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17655__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__B (.DIODE(_12244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17659__A (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17660__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17660__S (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17662__A (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17664__A (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17665__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17666__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17667__A (.DIODE(_12183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17668__A (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17669__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17670__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17670__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17671__A (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17675__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17676__A (.DIODE(_02861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17677__A (.DIODE(_12196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17678__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17679__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17679__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17683__A (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17684__A (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17685__A (.DIODE(_12204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17686__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17687__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17687__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17691__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17692__A (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17693__A (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17694__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17695__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17695__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17699__A (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17700__A (.DIODE(_02882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17701__A (.DIODE(_12220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17702__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17703__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17703__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17707__A (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17708__A (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17709__A (.DIODE(_12228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17710__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17715__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17716__A (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17717__A (.DIODE(_12236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17718__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17719__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17719__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17723__A (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17724__A (.DIODE(_02903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17725__A (.DIODE(_12244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17726__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17727__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17727__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17730__A (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17732__A (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17733__A (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17734__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17734__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17738__A (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17739__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__B1 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17744__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17745__A (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17746__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17747__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17751__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17752__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17753__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17757__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17758__A (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17759__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__A (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__A (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17765__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17769__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17770__A (.DIODE(_02942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17771__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17775__A (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17776__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17777__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17780__A (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17781__A (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17782__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17785__A (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17786__A (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17787__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17790__A (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17791__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17792__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17795__A (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17796__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17797__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17800__A (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17801__A (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17802__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17805__A (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17806__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17807__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17810__A (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17811__A (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17812__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17815__A (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17816__A (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17817__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17820__A (.DIODE(_12293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17821__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17822__A (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17823__A1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17823__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17824__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17826__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17828__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17830__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17832__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17834__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17836__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17838__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17843__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17844__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17848__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17849__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17852__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17853__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17854__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17857__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17858__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17862__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17865__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17866__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17869__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17870__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17873__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17874__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17878__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17881__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17884__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17887__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17890__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17893__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17896__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17902__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17905__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17908__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17909__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17909__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17912__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17912__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17918__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17918__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17921__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17921__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17927__A (.DIODE(_12292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17929__A (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__A1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17931__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17933__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17935__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17937__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17939__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17941__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17943__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17945__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17950__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17951__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17951__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17955__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17956__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17956__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17959__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17960__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17960__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17963__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17964__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17964__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17967__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17971__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17972__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17972__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17979__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17980__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17980__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17984__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17984__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17987__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17987__B1 (.DIODE(_03045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17990__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17994__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17997__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18000__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18003__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18006__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18012__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18015__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18018__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18021__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18024__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18027__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__A (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18035__A (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__A1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__A2 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18037__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18037__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18039__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18039__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18043__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18043__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18045__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18045__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18047__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18047__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__S (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18053__A (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18054__A (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18055__A (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18056__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18057__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18058__A (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18061__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18062__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18065__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18066__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18067__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18070__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18071__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18074__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18075__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18078__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18079__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18082__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18083__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18086__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18087__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18090__A (.DIODE(_03135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18091__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18094__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18097__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18100__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18103__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18106__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18109__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18112__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18115__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18118__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18121__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18122__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18125__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18125__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18134__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18134__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18141__A (.DIODE(_03207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18142__A (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18144__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18145__A1 (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18145__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18145__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18147__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18149__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18151__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18153__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18155__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18157__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18159__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18161__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18163__A (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18164__A (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__A (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18167__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18167__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18175__A (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18176__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18177__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18177__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18180__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18181__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18182__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18182__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18185__A (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18186__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18187__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18187__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18190__A (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18191__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18192__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18192__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18195__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18197__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18197__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18200__A (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18201__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__B1 (.DIODE(_12181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18205__A (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18206__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18207__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18211__A (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18212__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18215__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18216__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18219__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18220__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18223__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18224__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18227__A (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18228__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18231__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18232__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18235__A (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18236__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18239__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18242__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18245__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18248__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18251__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18257__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18260__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18263__A (.DIODE(_12293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18264__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18265__A1 (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18265__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18265__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18267__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18269__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18271__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18273__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18275__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18277__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18279__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18281__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18283__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18286__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18287__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18290__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18291__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18294__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18298__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18299__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18302__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18303__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18306__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18307__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18310__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18311__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18314__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18315__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18322__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18325__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18328__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18331__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18334__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18337__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18340__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18343__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18344__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18344__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18347__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18347__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18350__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18350__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18353__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18353__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18356__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18356__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18359__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18359__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18362__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18362__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18365__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18365__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18368__A (.DIODE(_12292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18369__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18370__A1 (.DIODE(_03372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18370__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18370__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18372__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18374__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18376__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18378__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18380__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18382__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18384__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18386__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18388__A (.DIODE(_03372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18389__A (.DIODE(_03372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18390__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18391__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18391__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18394__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18395__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18395__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18398__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18402__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18406__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18407__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18407__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18410__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18411__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18411__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18414__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18415__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18415__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18418__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18419__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18419__B1 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18422__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18423__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18430__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18433__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18436__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18439__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18442__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18445__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18448__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18451__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18454__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18457__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18460__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18463__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18469__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18472__A (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18473__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18474__A1 (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18474__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18474__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18476__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18478__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18480__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18486__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18488__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18490__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__A (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18494__A (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18495__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18496__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18499__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18503__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18504__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18507__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18508__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18511__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18512__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18515__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18516__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18519__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18520__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18523__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18524__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18527__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18529__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18531__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18532__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18534__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18535__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18537__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18538__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18540__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18541__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18543__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18544__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18546__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18547__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18549__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18550__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18552__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18556__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18557__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18559__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18560__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18562__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18563__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18565__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18566__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18568__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18569__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18571__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18572__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18574__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18575__S (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18578__A (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__A (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__B (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18581__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__A1 (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18586__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18586__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18588__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18588__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18590__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18590__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18592__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18592__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18594__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18594__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18598__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18598__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18600__A (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18601__A (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18602__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18603__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18604__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18606__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18607__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18608__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18610__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18611__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18612__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18614__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18618__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18619__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18620__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18622__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18624__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18626__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18627__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18628__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18630__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18631__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18632__S (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18634__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18639__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18642__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18645__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18648__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18651__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18654__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18657__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18660__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18663__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18666__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18669__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18672__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18675__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18678__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18681__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18684__A (.DIODE(_12293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18684__B (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18685__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__A1 (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18686__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18688__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18688__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18690__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18690__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18692__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18692__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18702__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18702__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18704__A (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18705__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18706__A (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18707__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18708__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18709__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18712__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18715__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18716__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18717__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18719__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18720__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18721__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18724__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18725__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18727__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18728__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18729__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18733__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18735__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18736__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18737__S (.DIODE(_03594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18739__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18743__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18744__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18747__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18750__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18752__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18753__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18755__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18756__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18758__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18759__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18761__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18762__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18764__A (.DIODE(_12180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18765__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18768__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18774__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18775__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18777__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18778__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18780__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18781__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18783__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18784__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18787__S (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18789__A (.DIODE(_12292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18789__B (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18790__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18791__A1 (.DIODE(_03665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18791__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18791__B1_N (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18793__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18793__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18795__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18795__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18797__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18797__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18799__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18799__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18801__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18801__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18803__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18803__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18805__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18805__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18807__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18807__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18809__A (.DIODE(_03665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18810__A (.DIODE(_03665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18811__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18812__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18813__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18815__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18816__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18817__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18819__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18820__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18821__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18823__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18824__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18825__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18827__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18828__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18829__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18831__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18832__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18833__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18835__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18836__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18837__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18839__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18840__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18841__S (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18843__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18844__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18845__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18849__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18852__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18855__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18858__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18861__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18864__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18867__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18876__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18879__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18882__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18885__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18888__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18894__A (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18894__B (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18895__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__A (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__A1 (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__A2 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18901__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18901__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18903__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18903__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18905__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18905__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18911__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18911__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18913__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18913__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18915__A (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18916__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18917__A (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18918__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18919__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18920__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18922__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18923__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18924__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18926__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18927__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18928__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18930__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18931__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18932__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18934__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18935__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18936__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18938__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18939__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18940__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18942__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18943__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18944__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18946__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18947__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__S (.DIODE(_03741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18954__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18960__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18963__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18966__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18969__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18972__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18975__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18976__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18976__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18979__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18979__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18982__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18982__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18985__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18985__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18988__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18988__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18991__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18991__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18994__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18994__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18997__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18997__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19000__A (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19000__B (.DIODE(_12175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19001__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19002__A (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__A1 (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19005__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19007__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19011__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19015__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19017__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19019__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19021__A (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19022__A (.DIODE(_03812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19023__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19024__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19024__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19027__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19028__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19028__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19031__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19035__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19036__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19036__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19039__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19040__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19040__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19043__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19044__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19044__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19047__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19048__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19048__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19051__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19052__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19052__B1 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19055__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19056__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19060__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19063__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19069__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19072__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19075__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19078__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19081__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19084__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19087__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19090__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19096__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19099__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19102__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__A (.DIODE(_12293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__B (.DIODE(_12175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19106__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19113__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19115__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19119__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19121__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19125__A (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19126__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19127__A (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19128__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19129__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19132__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19133__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19136__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19137__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19140__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19141__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19144__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19145__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19148__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19149__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19152__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19153__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19156__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19157__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19160__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19164__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19167__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19173__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19179__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19182__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19186__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19186__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19189__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19189__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19192__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19192__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19195__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19195__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19204__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19204__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19210__A (.DIODE(_12292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19210__B (.DIODE(_12175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19211__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19212__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19212__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19214__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19216__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19218__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19222__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19224__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19232__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19233__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19233__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19236__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19240__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19241__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19241__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19244__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19245__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19245__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19248__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19249__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19249__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19252__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19253__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19253__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19256__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19260__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__B1 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19264__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19265__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19269__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19272__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19275__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19278__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19281__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19284__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19287__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19290__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19293__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19296__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19299__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19302__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19305__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19308__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19311__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19314__B (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19315__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19315__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19317__A0 (.DIODE(_02810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19319__A0 (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19321__A0 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__A0 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19325__A0 (.DIODE(_02835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19327__A0 (.DIODE(_02839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19329__A0 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__A0 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19334__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19336__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19340__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19341__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19344__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19345__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19348__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19349__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19352__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19353__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19356__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19357__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19360__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19361__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19364__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19365__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19368__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19372__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19375__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19378__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19381__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19384__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19387__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19390__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19393__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19394__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19394__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19397__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19397__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19400__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19400__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19403__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19403__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19406__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19406__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19412__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19412__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19415__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19415__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19418__A (.DIODE(_02809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19420__C (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19421__B (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__A (.DIODE(_04103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19423__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19423__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19427__A (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19428__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19430__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19433__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19436__A (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19439__A (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19442__A (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19445__A (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19446__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19450__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19451__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19451__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19454__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19455__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19455__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19458__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19459__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19459__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19462__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19463__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19463__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19466__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19467__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19467__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19470__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19471__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19471__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19474__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19475__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19475__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19478__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19479__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19479__B1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19482__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19483__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19490__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19496__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19499__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19502__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19505__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19511__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19517__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19520__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19523__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19526__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19529__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19532__B (.DIODE(_12293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__A (.DIODE(_04103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19535__A1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19535__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19538__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19540__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19542__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19544__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19546__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19550__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19555__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19556__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19556__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19560__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19561__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19561__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19564__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19565__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19565__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19568__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19569__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19569__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19572__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19576__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19577__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19577__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19580__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19581__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19581__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19584__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19585__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19585__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19589__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19589__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19592__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19592__B1 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19595__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19596__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19596__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19599__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19599__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19602__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19602__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19605__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19605__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19608__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19608__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19611__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19611__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19614__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19614__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19617__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19617__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19620__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19620__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19623__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19623__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19626__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19626__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19629__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19629__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19632__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19632__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19635__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19635__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19638__B (.DIODE(_12292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19639__A (.DIODE(_04103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19639__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19641__A1 (.DIODE(_12290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19641__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19642__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19642__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19646__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19646__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19648__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19648__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19654__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19654__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19656__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19656__S (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19658__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19661__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19662__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19662__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19667__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19667__B1 (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19670__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19671__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19672__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19675__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19676__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19679__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19680__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19683__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19684__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19687__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19688__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19691__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19695__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19696__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19699__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19705__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19708__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19711__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19714__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19717__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19720__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19723__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19726__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19727__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19730__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19733__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19736__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19739__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19742__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19745__A (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__B (.DIODE(_12171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19747__A (.DIODE(_04103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19747__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19749__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19749__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19750__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19752__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19754__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19756__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19758__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19760__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19762__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19764__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19769__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19770__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19774__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19775__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19778__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19779__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19782__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19783__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19786__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19787__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19790__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19791__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19795__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19798__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19799__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19803__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19806__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19809__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19810__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19810__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19813__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19813__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19816__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19816__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19828__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19828__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19831__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19831__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19834__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19834__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19837__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19837__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19840__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19840__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19843__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19843__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19846__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19846__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19849__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19849__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__A (.DIODE(_03207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__C (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__A (.DIODE(_04407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19856__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19858__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19858__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19860__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19860__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19862__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19862__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19864__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19864__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19868__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19868__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19870__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19870__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19873__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19875__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19876__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19877__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19879__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19880__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19881__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19883__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19885__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19887__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19888__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19891__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19892__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19893__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19895__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19897__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19899__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19901__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19903__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19904__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19907__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19911__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19914__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19917__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19920__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19923__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19926__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19929__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19932__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19936__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19939__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19942__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19945__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19948__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19957__A (.DIODE(_04407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19957__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19959__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19960__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19962__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19964__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19966__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19968__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19970__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19979__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19980__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19980__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19984__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19985__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19985__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19988__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19989__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19990__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19993__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19994__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19997__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19998__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20001__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20002__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20005__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20006__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20009__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20010__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20014__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20017__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20020__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20023__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20029__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20032__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20035__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20038__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20041__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20044__A (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20048__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20048__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20051__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20051__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20054__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20054__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20057__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20057__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20060__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20060__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20063__A (.DIODE(_04407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20063__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20065__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20065__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20066__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20066__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20068__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20068__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20070__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20070__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20072__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20072__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20074__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20074__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20076__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20076__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20078__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20078__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20080__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20080__S (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20082__A (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20085__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20086__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20086__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20087__A (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20090__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20091__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20091__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20094__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20095__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20095__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20098__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20102__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20103__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20103__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20106__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20110__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20111__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20111__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20114__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20115__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20115__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20118__A (.DIODE(_04556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20119__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20119__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20122__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20122__B1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20125__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20126__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20127__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20133__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20139__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20142__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20148__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20151__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20154__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20157__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20160__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20163__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20166__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__A (.DIODE(_04407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20171__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20171__B1 (.DIODE(_02818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20172__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20174__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20176__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20178__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20180__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20182__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20184__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20186__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20191__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20192__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20196__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20197__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20200__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20201__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20202__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20205__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20206__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20209__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20210__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20213__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20214__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20217__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20218__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20221__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20222__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20226__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20229__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20232__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20235__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20238__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20241__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20244__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20247__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20250__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20253__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20256__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20257__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20257__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20260__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20260__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20263__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20263__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20266__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20266__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20269__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20269__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20272__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20272__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20275__A (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20275__C (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20276__A (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20276__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20277__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20277__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20279__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20279__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20281__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20281__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20283__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20283__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20285__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20285__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20287__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20287__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20289__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20289__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20291__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20291__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20293__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20293__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20297__B (.DIODE(_12185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20298__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20299__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20301__B (.DIODE(_12198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20302__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20303__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20305__B (.DIODE(_12206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20306__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20307__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20309__B (.DIODE(_12214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20310__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20311__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20313__B (.DIODE(_12222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20314__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20315__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20317__B (.DIODE(_12230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20318__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20321__B (.DIODE(_12238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20322__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20323__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20325__B (.DIODE(_12246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20326__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20327__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20329__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20330__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20334__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20337__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20340__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20343__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20346__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20349__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20352__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20355__A1 (.DIODE(_12170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20358__A1 (.DIODE(_12195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20361__A1 (.DIODE(_12203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20364__A1 (.DIODE(_12211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20367__A1 (.DIODE(_12219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20370__A1 (.DIODE(_12227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20373__A1 (.DIODE(_12235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20376__A1 (.DIODE(_12243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20379__A (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20379__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20381__A (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20382__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20382__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20383__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20385__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20389__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20391__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20393__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20395__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20397__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20402__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20403__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20403__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20407__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20408__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20408__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20411__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20412__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20412__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20419__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20420__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20420__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20423__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20424__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20424__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20427__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20428__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20428__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20431__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20432__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20432__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20436__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20436__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20439__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20439__B1 (.DIODE(_04689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20442__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20443__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20443__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20446__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20446__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20449__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20449__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20452__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20452__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20455__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20455__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20458__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20458__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20461__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20461__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20464__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20464__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20467__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20467__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20470__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20470__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20473__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20473__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20476__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20476__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20479__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20479__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20482__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20482__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20485__A (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20485__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20487__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20487__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20488__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20490__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20492__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20494__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20496__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20498__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20500__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20502__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20507__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20512__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20513__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20513__B1 (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20516__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20517__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20518__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20521__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20522__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20525__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20526__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20529__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20530__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20533__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20534__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20537__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20538__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20542__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20545__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20548__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20551__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20554__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20557__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20560__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20563__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20566__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20569__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20572__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20573__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20576__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20579__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20582__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20585__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20588__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20591__A (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20591__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20593__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20593__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20594__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20594__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20596__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20596__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20598__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20598__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20600__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20600__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20602__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20602__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20606__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20606__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20608__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20608__S (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20610__A (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20613__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20614__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20615__A (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20618__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20619__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20622__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20623__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20626__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20627__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20630__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20631__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20634__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20635__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20638__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20639__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20642__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20643__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20646__A (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20647__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20650__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20653__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20654__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20654__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20657__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20657__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20660__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20660__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20663__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20663__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20666__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20666__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20672__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20672__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20675__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20675__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20678__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20678__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20681__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20681__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20684__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20684__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20687__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20687__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20690__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20690__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20693__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20693__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20696__C (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20697__A (.DIODE(_04995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20697__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20698__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20698__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20700__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20702__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20704__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20706__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20708__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20710__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20712__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20714__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20717__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20719__A (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20720__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20721__A1 (.DIODE(_03222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20724__A (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20725__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20726__A1 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20729__A (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20730__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20731__A1 (.DIODE(_03232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20734__A (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20735__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20736__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20739__A (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20740__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20741__A1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20744__A (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20745__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20746__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20749__A (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20750__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20751__A1 (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20754__A (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20755__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20756__A1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20759__A1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20763__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20766__A1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20769__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20772__A1 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20775__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20778__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20781__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20784__A (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20785__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20786__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20786__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20789__A (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20790__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20790__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20793__A (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20794__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20794__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20797__A (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20798__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20798__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20801__A (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20802__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20802__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20805__A (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20806__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20806__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20809__A (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20810__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20810__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20813__A (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20814__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20814__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20817__A (.DIODE(_04995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20817__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20818__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20818__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20820__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20822__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20824__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20826__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20828__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20830__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20832__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20834__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20836__A (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20839__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20840__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20840__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20843__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20844__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20848__A (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20849__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20850__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20850__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20853__A (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20854__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20855__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20855__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20858__A (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20859__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20860__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20860__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20863__A (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20864__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20865__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20865__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20868__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20869__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20870__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20870__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20873__A (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20874__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20875__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20875__B1 (.DIODE(_05060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20878__A (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20879__A (.DIODE(_03702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20880__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20884__A (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20885__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20888__A (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20889__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20892__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20893__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20896__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20897__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20900__A (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20901__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20904__A (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20905__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20908__A (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20909__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20912__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20915__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20918__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20921__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20924__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20927__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20930__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20933__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20936__A (.DIODE(_04995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20936__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20937__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20937__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20939__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20939__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20941__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20941__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20943__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20943__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20945__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20945__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20947__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20947__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20949__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20949__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20951__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20951__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20953__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20953__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20956__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20957__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20959__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20960__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20961__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20963__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20964__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20965__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20967__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20968__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20969__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20971__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20972__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20973__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20975__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20976__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20977__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20979__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20980__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20981__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20983__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20984__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20985__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20987__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20988__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20989__S (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20991__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20995__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20998__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21001__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21004__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21007__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21010__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21013__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21016__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21017__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21020__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21023__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21026__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21029__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21032__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21035__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21038__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21041__A (.DIODE(_04995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21041__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21044__A0 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21046__A0 (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21048__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21050__A0 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21052__A0 (.DIODE(_04115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21054__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21056__A0 (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21058__A0 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21063__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21064__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21064__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21068__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21069__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21069__B1 (.DIODE(_04966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21072__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21073__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21074__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21077__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21078__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21081__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21082__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21085__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21086__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21089__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21090__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21093__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21094__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21098__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21101__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21104__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21107__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21110__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21113__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21116__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21119__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21122__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21125__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21128__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21129__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21129__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21132__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21132__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21135__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21135__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21138__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21138__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21141__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21141__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21144__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21144__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21147__A (.DIODE(_02809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21149__A (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21149__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21150__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21150__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21152__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21154__A (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21157__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21158__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21160__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21161__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21163__A (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21164__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21166__A (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21167__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21169__A (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21170__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21172__A (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21173__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21177__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21178__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21181__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21182__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21185__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21186__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21189__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21190__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21193__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21194__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21197__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21198__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21201__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21202__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21205__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21206__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21209__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21210__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21214__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21217__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21220__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21223__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21226__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21229__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21232__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21235__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21238__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21241__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21244__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21247__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21250__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21253__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21256__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21259__A (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21259__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21261__A1 (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21261__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21262__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21264__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21266__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21268__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21270__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21272__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21274__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21276__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21281__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21282__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21282__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21286__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21287__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21287__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21290__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21291__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21291__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21294__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21295__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21295__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21298__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21299__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21299__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21302__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21303__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21303__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21306__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21307__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21307__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21310__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21311__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21311__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21318__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21318__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21321__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21322__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21322__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21325__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21325__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21328__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21328__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21331__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21331__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21334__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21334__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21337__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21337__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21340__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21340__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21343__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21343__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21346__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21346__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21349__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21349__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21352__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21352__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21355__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21355__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21358__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21358__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21361__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21361__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21364__A (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21365__A (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21365__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21367__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21367__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21368__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21368__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21370__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21370__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21372__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21372__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21374__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21374__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21376__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21376__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21378__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21378__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21380__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21380__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21382__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21382__S (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21384__A (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21385__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21388__A (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21389__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21389__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21390__A (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21393__A (.DIODE(_02861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21394__A (.DIODE(_02863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21395__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21395__B1 (.DIODE(_05442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21398__A (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21399__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21400__A (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21401__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21404__A (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21405__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21406__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21409__A (.DIODE(_02882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21410__A (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21411__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21414__A (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21415__A (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21416__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21419__A (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21420__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21421__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21424__A (.DIODE(_02903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21425__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21426__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21429__A (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21430__A (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21431__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21434__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21435__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21438__A (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21439__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21442__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21443__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21446__A (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21447__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21450__A (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21451__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21454__A (.DIODE(_02942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21455__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21458__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21459__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21462__A (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21463__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21466__A (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21467__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21470__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21471__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21472__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21475__A (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21476__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21479__A (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21480__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21483__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21484__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21487__A (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21488__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21491__A (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21492__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21495__A (.DIODE(_05319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21495__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21497__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21497__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21498__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21498__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21500__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21500__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21502__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21502__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21504__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21504__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21506__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21506__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21508__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21508__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21510__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21510__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21512__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21512__S (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21514__A (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21516__A (.DIODE(_12183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21518__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21519__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21520__A (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21523__A (.DIODE(_12196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21524__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21525__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21528__A (.DIODE(_12204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21529__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21530__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21533__A (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21534__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21535__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21538__A (.DIODE(_12220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21539__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21540__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21543__A (.DIODE(_12228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21544__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21545__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21548__A (.DIODE(_12236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21549__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21550__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21553__A (.DIODE(_12244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21554__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21555__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21558__A (.DIODE(_05572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21559__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21562__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21565__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21566__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21569__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21572__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21575__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21578__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21581__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21584__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21587__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21590__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21593__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21596__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21599__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21602__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21605__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21608__A (.DIODE(_03207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21609__A (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21609__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21610__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21610__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21612__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21614__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21616__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21618__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21620__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21622__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21624__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21626__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21629__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21631__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21632__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21635__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21636__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21639__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21640__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21643__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21644__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21647__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21648__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21651__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21652__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21655__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21656__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21659__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21660__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21663__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21667__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21670__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21673__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21676__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21679__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21682__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21685__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21688__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21689__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21689__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21692__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21692__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21695__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21695__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21698__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21698__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21701__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21701__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21704__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21704__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21707__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21707__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21710__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21710__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21713__A (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21713__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21715__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21715__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21716__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21718__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21720__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21722__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21724__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21726__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21728__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21730__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21735__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21736__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21740__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21741__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21744__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21745__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21746__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21749__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21750__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21753__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21754__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21757__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21758__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21761__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21762__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21765__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21766__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21770__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21773__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21776__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21779__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21782__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21785__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21788__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21791__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21794__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21797__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21800__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21801__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21801__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21804__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21804__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21807__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21807__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21810__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21810__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21813__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21813__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21816__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21816__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21819__A (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21819__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21821__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21821__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21822__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21822__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21824__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21824__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21826__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21826__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21828__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21828__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21830__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21830__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21832__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21832__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21834__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21834__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21836__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21836__S (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21838__A (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21841__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21842__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21842__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21843__A (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21846__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21847__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21847__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21850__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21851__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21851__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21854__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21855__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21855__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21858__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21859__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21859__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21862__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21863__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21863__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21866__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21867__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21867__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21870__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21871__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21871__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21874__A (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21875__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21875__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21878__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21878__B1 (.DIODE(_05785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21881__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21882__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21885__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21888__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21891__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21894__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21897__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21900__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21903__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21906__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21909__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21912__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21915__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21918__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21921__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21924__A (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21924__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21926__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21926__B1 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21927__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21929__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21931__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21933__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21935__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21937__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21939__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21941__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21946__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21947__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21951__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21952__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21955__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21956__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21957__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21958__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21961__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21962__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21965__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21966__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21969__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21970__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21973__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21974__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21977__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21978__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21982__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21985__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21988__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21991__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21994__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21997__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22000__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22003__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22006__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22009__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22012__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22013__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22013__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22016__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22016__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22019__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22019__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22022__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22022__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22025__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22025__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22028__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22028__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22031__A (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22032__A (.DIODE(_05946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22032__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22033__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22033__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22035__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22035__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22037__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22037__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22039__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22039__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22041__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22041__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22043__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22043__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22045__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22045__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22047__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22047__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22049__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22049__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22053__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22054__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22054__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22055__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22057__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22058__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22058__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22059__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22061__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22062__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22062__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22063__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22065__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22066__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22066__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22067__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22069__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22070__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22070__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22071__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22073__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22074__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22074__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22075__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22077__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22078__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22078__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22079__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22081__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22082__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22082__B1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22083__S (.DIODE(_05949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22085__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22086__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22090__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22093__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22096__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22099__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22102__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22105__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22108__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22111__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22114__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22117__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22120__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22123__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22126__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22129__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22132__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22135__A (.DIODE(_05946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22135__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22137__A (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22138__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22138__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22139__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22139__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22141__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22141__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22143__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22143__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22145__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22145__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22147__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22147__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22149__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22149__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22151__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22151__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22153__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22153__S (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22155__A (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22158__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22159__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22159__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22160__A (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22163__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22164__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22164__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22167__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22168__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22168__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22171__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22172__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22172__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22175__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22176__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22176__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22179__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22180__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22180__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22183__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22184__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22184__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22187__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22188__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22188__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22191__A (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22192__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22192__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22195__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22195__B1 (.DIODE(_05933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22198__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22199__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22202__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22205__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22208__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22211__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22214__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22217__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22220__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22223__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22226__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22229__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22232__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22235__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22238__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22241__A (.DIODE(_05946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22241__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22243__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22243__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22244__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22246__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22248__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22250__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22252__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22254__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22256__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22258__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22263__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22264__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22268__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22269__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22272__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22273__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22274__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22277__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22278__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22281__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22282__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22285__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22286__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22289__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22290__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22293__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22294__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22298__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22301__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22304__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22307__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22310__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22313__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22316__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22319__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22322__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22325__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22328__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22329__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22332__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22335__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22338__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22341__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22344__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22347__A (.DIODE(_05946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22347__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22349__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22349__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22350__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22350__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22352__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22352__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22354__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22354__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22356__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22356__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22358__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22358__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22360__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22360__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22362__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22362__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22364__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22364__S (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22366__A (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22369__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22370__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22371__A (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22374__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22375__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22378__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22379__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22382__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22383__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22386__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22387__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22390__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22391__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22394__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22395__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22398__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22399__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22402__A (.DIODE(_06168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22403__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22406__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22409__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22410__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22410__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22413__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22413__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22416__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22416__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22419__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22419__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22422__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22422__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22425__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22425__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22428__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22428__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22431__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22431__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22434__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22434__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22437__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22437__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22440__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22440__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22443__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22443__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22446__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22446__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22449__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22449__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22453__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22453__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22454__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22454__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22456__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22458__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22460__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22462__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22464__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22466__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22468__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22470__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22473__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22475__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22476__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22479__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22480__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22483__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22484__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22487__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22488__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22491__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22492__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22495__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22496__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22499__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22500__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22503__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22504__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22507__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22511__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22514__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22517__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22520__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22523__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22526__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22529__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22532__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22533__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22533__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22536__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22536__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22539__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22539__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22542__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22542__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22545__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22545__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22548__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22548__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22551__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22551__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22554__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22554__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22557__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22557__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22558__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22558__B1_N (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22560__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22562__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22564__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22566__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22568__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22570__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22572__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22574__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22578__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22579__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22579__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22582__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22583__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22583__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22586__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22587__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22587__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22590__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22591__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22591__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22594__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22595__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22595__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22598__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22599__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22599__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22602__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22603__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22603__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22606__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22607__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22607__B1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22610__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22611__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22615__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22618__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22621__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22624__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22627__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22630__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22633__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22636__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22639__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22642__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22645__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22648__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22651__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22654__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22657__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22660__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22660__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22661__A (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22662__A2 (.DIODE(_03813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22662__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22664__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22664__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22666__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22666__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22668__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22668__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22670__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22670__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22672__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22672__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22674__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22674__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22676__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22676__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22678__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22678__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22681__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22683__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22684__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22685__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22687__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22688__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22689__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22691__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22692__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22693__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22695__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22696__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22697__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22699__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22700__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22701__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22703__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22704__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22705__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22707__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22708__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22709__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22711__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22712__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22713__S (.DIODE(_06386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22715__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22719__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22722__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22725__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22728__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22731__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22734__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22737__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22740__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22741__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22741__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22744__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22744__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22747__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22747__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22750__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22750__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22753__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22753__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22756__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22756__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22759__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22759__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22762__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22762__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22765__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22765__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22767__A1 (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22767__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22768__A0 (.DIODE(_05318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22770__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22772__A0 (.DIODE(_05326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22774__A0 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22776__A0 (.DIODE(_05330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22778__A0 (.DIODE(_05332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22780__A0 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22782__A0 (.DIODE(_05336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22787__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22788__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22788__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22792__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22793__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22793__B1 (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22796__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22797__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22798__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22801__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22802__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22805__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22806__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22809__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22810__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22813__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22814__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22817__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22818__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22822__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22825__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22828__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22831__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22834__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22837__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22840__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22843__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22846__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22849__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22852__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22853__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22853__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22856__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22856__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22859__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22859__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22862__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22862__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22865__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22865__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22868__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22868__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22871__A (.DIODE(_02809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22874__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22874__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22875__A (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22876__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22876__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22878__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22880__A (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22881__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22883__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22884__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22886__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22887__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22889__A (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22890__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22892__A (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22893__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22895__A (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22896__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22898__A (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22899__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22903__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22904__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22904__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22907__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22908__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22908__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22911__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22912__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22912__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22915__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22916__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22916__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22919__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22920__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22920__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22923__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22924__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22924__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22927__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22928__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22928__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22931__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22932__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22932__B1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22935__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22936__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22940__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22943__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22946__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22949__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22952__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22955__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22958__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22961__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22964__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22967__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22970__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22973__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22976__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22979__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22982__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22985__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22985__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22986__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22986__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22988__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22990__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22992__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22994__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22996__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22998__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23000__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23002__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23005__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23007__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23008__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23011__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23012__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23015__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23016__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23019__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23020__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23023__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23024__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23027__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23028__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23031__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23032__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23035__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23036__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23039__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23043__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23046__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23049__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23052__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23055__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23058__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23061__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23064__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23065__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23068__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23071__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23074__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23077__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23080__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23083__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23086__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23089__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23089__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23090__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23090__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23092__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23094__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23096__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23098__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23100__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23102__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23104__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23106__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23110__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23111__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23114__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23115__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23118__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23119__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23122__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23123__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23126__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23127__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23130__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23131__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23134__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23135__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23138__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23139__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23142__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23143__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23145__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23147__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23148__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23150__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23151__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23153__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23154__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23156__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23157__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23159__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23160__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23162__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23163__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23165__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23166__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23168__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23169__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23171__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23172__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23174__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23175__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23177__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23178__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23180__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23181__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23183__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23184__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23186__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23187__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23189__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23190__S (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23192__A (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23193__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23193__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23195__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23195__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23196__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23196__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23198__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23198__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23200__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23200__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23202__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23202__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23204__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23204__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23206__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23206__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23208__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23208__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23210__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23210__S (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23212__A (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23215__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23216__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23216__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23217__A (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23220__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23221__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23221__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23224__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23225__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23225__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23228__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23229__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23229__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23232__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23233__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23233__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23236__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23237__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23237__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23240__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23241__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23241__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23244__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23245__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23245__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23248__A (.DIODE(_06758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23249__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23249__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23252__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23252__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23255__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23256__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23259__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23262__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23265__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23268__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23271__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23274__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23277__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23280__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23283__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23286__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23289__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23292__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23295__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23298__A (.DIODE(_03207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23299__A (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23299__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23300__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23300__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23302__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23302__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23304__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23304__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23306__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23306__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23308__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23308__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23310__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23310__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23312__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23312__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23314__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23314__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23316__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23316__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23319__A (.DIODE(_05183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23321__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23322__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23323__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23325__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23326__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23327__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23329__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23330__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23331__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23333__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23334__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23335__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23337__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23338__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23339__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23341__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23342__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23343__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23345__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23346__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23347__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23349__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23350__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23351__S (.DIODE(_06832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23353__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23357__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23360__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23363__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23366__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23369__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23372__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23375__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23378__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__23379__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23380__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23383__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23386__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23389__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23392__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23395__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23398__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23401__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23404__A (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23404__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23405__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23405__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23407__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23409__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23411__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23413__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23415__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23417__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23419__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23421__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23425__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23426__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23429__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23430__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23433__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23434__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23437__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23438__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23441__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23442__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23445__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23446__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23449__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23450__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23453__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23454__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23457__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23458__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23462__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23465__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23468__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23471__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23474__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23477__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23480__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23483__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23486__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23489__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23492__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23495__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23498__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23501__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23504__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23507__A (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23507__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23508__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23508__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23510__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23512__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23514__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23516__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23518__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23520__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23522__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23524__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23527__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23529__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23530__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23533__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23534__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23537__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23538__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23541__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23542__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23545__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23546__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23549__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23550__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23553__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23554__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23557__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23558__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23561__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23565__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23568__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23571__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23574__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23577__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23580__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23583__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23586__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23587__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23587__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23590__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23590__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23593__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23593__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23596__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23596__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23599__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23599__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23602__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23602__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23605__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23605__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23608__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23608__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23611__A (.DIODE(_06829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23611__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23613__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23613__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23614__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23616__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23618__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23620__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23622__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23624__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23626__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23628__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23633__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23634__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23638__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23639__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23642__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23643__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23644__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23647__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23648__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23651__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23652__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23655__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23656__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23659__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23660__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23663__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23664__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23668__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23671__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23674__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23677__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23680__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23683__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23686__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23689__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23692__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23695__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23698__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23699__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23699__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23702__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23702__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23705__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23705__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23708__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23708__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23711__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23711__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23714__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23714__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23717__A (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23718__B (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23719__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23719__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23721__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23721__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23723__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23723__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23725__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23725__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23727__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23727__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23729__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23729__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23731__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23731__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23733__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23733__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23735__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23735__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23739__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23740__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23740__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23741__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23743__B (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23744__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23744__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23745__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23747__B (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23748__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23748__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23749__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23751__B (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23752__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23752__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23753__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23755__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23756__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23756__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23757__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23759__B (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23760__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23760__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23761__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23763__B (.DIODE(_05034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23764__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23764__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23765__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23767__B (.DIODE(_05038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23768__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23768__B1 (.DIODE(_07029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23769__S (.DIODE(_07123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23771__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23772__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23776__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23779__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23782__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23785__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23788__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23791__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23794__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23797__A1 (.DIODE(_05059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23800__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23803__A1 (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23806__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23809__A1 (.DIODE(_05072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23812__A1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23815__A1 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23818__A1 (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23821__B (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23822__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23822__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23824__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23826__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23828__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23830__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23832__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23834__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23836__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23838__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23841__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23843__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23844__A1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23847__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23848__A1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23851__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23852__A1 (.DIODE(_05105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23855__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23856__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23859__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23860__A1 (.DIODE(_05113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23863__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23864__A1 (.DIODE(_05117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23867__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23868__A1 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23871__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23872__A1 (.DIODE(_05125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23875__A1 (.DIODE(_05129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23879__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23882__A1 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23885__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23888__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23891__A1 (.DIODE(_05146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23894__A1 (.DIODE(_05149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23897__A1 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23900__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23901__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23904__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23907__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23910__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23913__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23916__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23919__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23922__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23925__B (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23926__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23926__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23928__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23930__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23932__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23934__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23936__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23938__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23940__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23942__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23946__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23947__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23950__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23951__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23954__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23955__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23958__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23959__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23962__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23963__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23966__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23967__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23970__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23971__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23974__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23975__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23978__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23979__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23983__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23986__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23989__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23992__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23995__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23998__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24001__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24004__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24007__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24010__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24013__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24016__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24019__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24022__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24025__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24028__B (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24030__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24030__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24031__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24033__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24035__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24037__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24039__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24041__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24043__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24045__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24050__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24051__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24051__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24055__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24056__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24056__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24059__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24060__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24060__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24063__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24064__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24064__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24067__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24068__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24068__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24071__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24072__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24072__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24075__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24076__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24076__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24079__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24080__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24080__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24084__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24084__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24087__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24087__B1 (.DIODE(_07107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24090__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24091__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24091__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24094__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24094__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24097__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24097__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24100__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24100__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24103__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24103__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24106__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24106__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24109__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24109__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24112__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24112__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24115__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24115__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24118__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24118__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24121__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24121__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24124__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24124__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24127__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24127__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24130__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24130__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24133__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24133__B (.DIODE(_12311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24135__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24135__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24136__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24138__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24140__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24142__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24144__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24146__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24148__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24150__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24155__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24156__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24156__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24160__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24161__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24161__B1 (.DIODE(_07379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24164__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24165__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24166__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24169__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24170__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24173__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24174__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24177__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24178__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24181__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24182__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24185__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24186__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24190__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24193__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24196__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24199__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24202__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24205__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24208__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24211__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24214__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24217__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24220__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24221__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24224__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24227__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24230__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24233__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24236__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24239__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24239__B (.DIODE(_12311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24241__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24241__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24242__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24244__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24246__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24248__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24250__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24252__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24254__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24256__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24261__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24262__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24266__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24267__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24270__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24271__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24274__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24275__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24278__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24279__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24282__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24283__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24286__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24287__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24290__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24291__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24295__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24298__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24301__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24302__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24305__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24308__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24311__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24314__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24317__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24320__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24323__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24326__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24329__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24332__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24335__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24338__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24341__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24344__A (.DIODE(_04257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24344__B (.DIODE(_12311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24346__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24346__B1 (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24347__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24349__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24351__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24353__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24355__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24357__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24359__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24361__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24366__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24367__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24371__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24372__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24375__A (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24376__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24377__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24380__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24381__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24384__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24385__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24388__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24389__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24392__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24393__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24396__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24397__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24401__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24404__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24407__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24410__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24413__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24416__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24419__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24422__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24425__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24428__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24431__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24432__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24432__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24435__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24435__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24438__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24438__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24441__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24441__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24444__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24444__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24447__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24447__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24451__A (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24452__A1 (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24452__B1 (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24454__A0 (.DIODE(_06530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24456__A0 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24458__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24460__A0 (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24462__A0 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24464__A0 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24466__A0 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24468__A0 (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24471__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24471__A2 (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24471__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24472__A1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24475__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24475__A2 (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24475__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24476__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24479__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24479__A2 (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24479__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24480__A1 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24483__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24483__A2 (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24483__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24484__A1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24487__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24487__A2 (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24487__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24488__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24491__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24491__A2 (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24491__B1 (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24492__A1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24495__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24495__A2 (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24495__B1 (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24496__A1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24499__A1 (.DIODE(_07629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24499__A2 (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24499__B1 (.DIODE(_09129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24500__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24503__A1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24505__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24507__A1 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24508__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24510__A1 (.DIODE(_02922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24511__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24513__A1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24514__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24516__A1 (.DIODE(_02933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24517__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24519__A1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24520__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24522__A1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24523__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24525__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24526__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24528__A1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24529__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24531__A1 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24532__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24534__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24535__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24537__A1 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24538__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24540__A1 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24541__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24543__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24544__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24546__A1 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24547__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24549__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24550__S (.DIODE(_07667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24552__A (.DIODE(_02809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24553__A (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24554__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24554__B1 (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24555__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24555__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24557__A (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24558__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24558__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24560__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24561__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24561__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24563__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24564__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24564__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24566__A (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24567__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24567__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24569__A (.DIODE(_02838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24570__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24570__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24572__A (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24573__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24573__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24575__A (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24576__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24576__S (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24578__A (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24581__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24582__A1 (.DIODE(_05484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24582__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24583__A (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24586__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24587__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24587__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24590__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24591__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24591__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24594__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24595__A1 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24595__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24598__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24599__A1 (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24599__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24602__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24603__A1 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24603__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24606__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24607__A1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24607__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24610__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24611__A1 (.DIODE(_05516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24611__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24614__A (.DIODE(_07701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24615__A1 (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24615__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24618__A1 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24618__B1 (.DIODE(_07616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24621__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24622__A1 (.DIODE(_05527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24625__A1 (.DIODE(_05530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24628__A1 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24631__A1 (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24634__A1 (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24637__A1 (.DIODE(_05542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24640__A1 (.DIODE(_05545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24643__A1 (.DIODE(_05548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24646__A1 (.DIODE(_05551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24649__A1 (.DIODE(_05555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24652__A1 (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24655__A1 (.DIODE(_05561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24658__A1 (.DIODE(_05564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24661__A1 (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24664__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24666__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24666__B1 (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24667__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24669__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24671__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24673__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24675__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24677__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24679__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24681__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24686__A (.DIODE(_05583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24687__A1 (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24691__A (.DIODE(_05589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24692__A1 (.DIODE(_02861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24695__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24696__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24697__A1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24700__A (.DIODE(_05597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24701__A1 (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24704__A (.DIODE(_05601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24705__A1 (.DIODE(_02882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24708__A (.DIODE(_05605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24709__A1 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24712__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24713__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24716__A (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24717__A1 (.DIODE(_02903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24721__A1 (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24724__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24727__A1 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24730__A1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24733__A1 (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24736__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24739__A1 (.DIODE(_02942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24742__A1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24745__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24748__A1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24751__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24752__A1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24752__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24755__A1 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24755__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24758__A1 (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24758__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24761__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24761__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24764__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24764__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24767__A1 (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24767__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24772__A1 (.DIODE(_06755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24772__B1 (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24773__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24773__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24775__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24775__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24777__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24777__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24779__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24779__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24781__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24781__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24783__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24783__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24785__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24785__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24787__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24787__S (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24789__A (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24792__A (.DIODE(_12183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24793__A1 (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24793__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24794__A (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24797__A (.DIODE(_12196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24798__A1 (.DIODE(_02861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24798__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24801__A (.DIODE(_12204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24802__A1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24802__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24805__A (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24806__A1 (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24806__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24809__A (.DIODE(_12220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24810__A1 (.DIODE(_02882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24810__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24813__A (.DIODE(_12228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24814__A1 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24814__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24817__A (.DIODE(_12236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24818__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24818__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24821__A (.DIODE(_12244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24822__A1 (.DIODE(_02903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24822__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24825__A (.DIODE(_07855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24826__A1 (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24826__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24829__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24829__B1 (.DIODE(_07840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24832__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24833__A1 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24833__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24836__A1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24836__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24839__A1 (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24839__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24842__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24842__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24845__A1 (.DIODE(_02942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24845__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24848__A1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24848__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24851__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24851__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24854__A1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24854__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24857__A1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24857__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24860__A1 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24860__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24863__A1 (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24863__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24866__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24866__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24869__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24869__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24872__A1 (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24872__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24875__A (.DIODE(_12313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24876__A1 (.DIODE(_12289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24876__B1 (.DIODE(_12190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24877__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24877__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24879__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24879__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24881__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24881__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24883__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24883__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24885__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24885__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24887__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24887__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24889__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24889__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24891__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24891__S (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24893__A (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24896__A (.DIODE(_12183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24897__A1 (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24897__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24898__A (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24901__A (.DIODE(_12196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24902__A1 (.DIODE(_02861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24902__B1 (.DIODE(_07897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24905__A (.DIODE(_09057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24906__A (.DIODE(_12204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24907__A1 (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24910__A (.DIODE(_12212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24911__A1 (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24914__A (.DIODE(_12220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24915__A1 (.DIODE(_02882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24918__A (.DIODE(_12228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24919__A1 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24922__A (.DIODE(_12236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24923__A1 (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24926__A (.DIODE(_12244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24927__A1 (.DIODE(_02903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24930__A (.DIODE(_07927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24931__A1 (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24934__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24937__A1 (.DIODE(_02921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24940__A1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24943__A1 (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24946__A1 (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24949__A1 (.DIODE(_02942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24952__A1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24955__A1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24958__A1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24961__A1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24961__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24964__A1 (.DIODE(_02963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24964__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24967__A1 (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24967__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24970__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24970__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24973__A1 (.DIODE(_02975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24973__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24976__A1 (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24976__B1 (.DIODE(_12851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24979__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24980__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24980__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24982__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24984__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24986__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24988__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24990__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24992__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24994__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24996__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24999__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25001__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25002__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25005__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25006__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25009__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25010__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25013__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25014__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25017__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25018__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25021__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25022__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25025__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25026__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25029__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25030__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25033__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25037__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25040__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25043__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25046__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25049__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25052__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25055__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25058__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25059__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25059__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25062__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25062__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25065__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25065__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25068__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25068__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25071__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25071__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25074__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25074__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25077__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25077__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25080__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25080__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25083__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25084__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25084__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25086__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25086__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25088__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25088__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25090__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25090__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25092__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25092__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25094__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25094__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25096__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25096__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25098__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25098__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25100__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25100__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25104__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25105__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25105__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25106__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25108__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25109__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25109__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25110__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25112__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25113__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25113__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25114__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25116__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25117__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25117__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25118__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25120__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25121__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25121__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25122__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25124__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25125__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25125__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25126__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25128__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25129__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25129__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25130__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25132__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25133__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25133__B1 (.DIODE(_08053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25134__S (.DIODE(_08072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25136__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25137__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25141__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25144__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25147__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25150__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25153__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25156__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25159__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25162__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25165__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25168__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25171__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25174__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25177__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25180__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25183__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25186__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25187__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25187__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25189__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25191__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25193__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25195__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25197__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25199__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25201__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25203__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25206__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25208__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25209__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25212__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25213__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25216__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25217__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25220__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25221__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25224__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25225__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25228__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25229__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25232__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25233__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25236__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25237__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25240__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25244__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25247__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25250__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25253__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25256__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25259__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25262__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25265__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25266__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25266__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25269__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25269__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25272__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25272__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25275__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25275__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25278__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25278__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25281__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25281__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25284__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25284__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25287__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25287__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25290__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25291__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25291__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25293__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25295__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25297__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25299__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25301__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25303__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25305__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25307__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25311__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25312__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25312__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25315__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25316__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25316__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25319__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25320__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25320__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25323__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25324__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25324__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25327__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25328__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25328__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25331__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25332__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25332__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25335__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25336__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25336__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25339__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25340__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25340__B1 (.DIODE(_08196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25343__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25344__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25348__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25351__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25354__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25357__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25360__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25363__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25366__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25369__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25372__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25375__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25378__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25381__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25384__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25387__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25390__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25393__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25394__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25394__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25396__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25396__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25398__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25398__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25400__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25400__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25402__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25402__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25404__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25404__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25406__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25406__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25408__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25408__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25410__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25410__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25413__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25415__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25416__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25417__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25419__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25420__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25421__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25423__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25424__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25425__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25427__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25428__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25429__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25431__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25432__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25433__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25435__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25436__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25437__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25439__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25440__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25441__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25443__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25444__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25445__S (.DIODE(_08286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25447__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25451__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25454__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25457__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25460__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25463__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25466__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25469__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25472__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25473__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25476__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25479__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25482__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25485__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25488__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25491__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25494__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25497__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25498__A1 (.DIODE(_08356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25498__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25498__B1_N (.DIODE(_06384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25500__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25502__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25504__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25506__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25508__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25510__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25512__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25514__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25516__A (.DIODE(_08356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25517__A (.DIODE(_08356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25518__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25519__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25522__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25523__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25526__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25527__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25530__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25531__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25534__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25535__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25538__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25539__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25542__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25543__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25546__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25547__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25550__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25551__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25555__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25558__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25561__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25564__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25567__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25570__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25573__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25576__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25579__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25582__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25585__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25588__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25591__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25594__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25597__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25600__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25601__A2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25601__B1_N (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25603__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25605__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25607__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25609__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25611__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25613__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25615__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25617__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25620__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25622__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25623__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25626__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25627__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25630__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25631__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25634__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25635__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25638__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25639__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25642__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25643__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25646__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25647__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25650__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25651__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25654__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25658__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25661__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25664__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25667__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25670__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25673__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25676__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25679__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25680__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25680__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25683__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25683__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25686__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25686__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25689__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25689__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25692__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25692__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25695__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25695__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25698__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25698__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25701__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25701__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25704__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25705__A2 (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25705__B1_N (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25707__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25709__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25711__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25713__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25715__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25717__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25719__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25721__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25725__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25726__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25726__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25729__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25730__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25730__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25733__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25734__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25734__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25737__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25738__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25738__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25741__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25742__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25742__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25745__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25746__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25746__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25749__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25750__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25750__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25753__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25754__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25754__B1 (.DIODE(_08482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25757__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25758__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25762__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25765__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25768__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25771__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25774__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25777__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25780__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25783__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25786__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25789__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25792__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25795__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25798__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25801__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25804__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25807__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25808__A2 (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25808__B1_N (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25810__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25810__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25812__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25812__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25814__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25814__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25816__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25816__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25818__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25818__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25820__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25820__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25822__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25822__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25824__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25824__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25827__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25829__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25830__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25831__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25833__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25834__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25835__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25837__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25838__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25839__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25841__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25842__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25843__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25845__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25846__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25847__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25849__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25850__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25851__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25853__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25854__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25855__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25857__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25858__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25859__S (.DIODE(_08572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25861__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25865__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25868__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25871__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25874__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25877__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25880__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25883__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25886__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25887__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25887__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25890__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25890__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25893__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25893__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25896__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25896__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25899__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25899__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25902__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25902__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25905__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25905__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25908__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25908__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25911__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25912__A2 (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25912__B1_N (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25914__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25916__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25918__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25920__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25922__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25924__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25926__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25928__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25932__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25933__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25933__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25936__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25937__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25937__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25940__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25941__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25941__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25944__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25945__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25945__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25948__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25949__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25949__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25952__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25953__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25953__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25956__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25957__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25957__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25960__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25961__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25961__B1 (.DIODE(_08625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25964__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25965__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25969__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25972__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25975__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25978__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25981__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25984__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25987__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25990__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25993__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25996__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25999__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26002__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26005__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26008__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26011__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26014__B (.DIODE(_12177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26015__A2 (.DIODE(_09109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26015__B1_N (.DIODE(_12189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26017__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26017__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26019__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26019__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26021__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26021__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26023__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26023__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26025__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26025__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26027__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26027__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26029__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26029__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26031__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26031__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26034__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26036__B (.DIODE(_12184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26037__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26038__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26040__B (.DIODE(_12197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26041__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26042__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26044__B (.DIODE(_12205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26045__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26046__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26048__B (.DIODE(_12213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26049__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26050__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26052__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26053__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26054__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26056__B (.DIODE(_12229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26057__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26058__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26060__B (.DIODE(_12237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26061__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26062__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26064__B (.DIODE(_12245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26065__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26066__S (.DIODE(_08715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26068__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26072__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26075__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26078__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26081__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26084__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26087__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26090__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26093__A (.DIODE(_09125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26094__A1 (.DIODE(_12169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26094__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26097__A1 (.DIODE(_12194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26097__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26100__A1 (.DIODE(_12202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26100__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26103__A1 (.DIODE(_12210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26103__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26106__A1 (.DIODE(_12218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26106__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26109__A1 (.DIODE(_12226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26109__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26112__A1 (.DIODE(_12234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26112__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26115__A1 (.DIODE(_12242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26115__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26118__A0 (.DIODE(_07699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26118__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26120__A0 (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26120__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26122__A0 (.DIODE(_07705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26122__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26124__A0 (.DIODE(_07707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26124__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26126__A0 (.DIODE(_07709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26126__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26128__A0 (.DIODE(_07711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26128__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26130__A0 (.DIODE(_07713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26130__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26132__A0 (.DIODE(_07715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26132__S (.DIODE(_12192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26134__A1 (.DIODE(_02850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26134__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26138__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26138__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26141__A1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26141__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26144__A1 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26144__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26147__A1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26147__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26150__A1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26150__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26153__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26153__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26156__A1 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26156__B1 (.DIODE(_08768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26159__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26159__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26162__A1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26162__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26165__A1 (.DIODE(_02920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26165__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26168__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26168__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26171__A1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26171__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26174__A1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26174__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26177__A1 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26177__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26180__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26180__B1 (.DIODE(_12840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26183__B_N (.DIODE(_09128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26185__A2 (.DIODE(_09105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26185__B1 (.DIODE(_12328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26186__A0 (.DIODE(_09107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26199__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26200__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26201__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26202__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26203__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26204__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26205__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26206__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26213__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26214__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26253__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26254__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26255__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26263__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26264__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26265__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26266__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26268__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26269__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26270__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26271__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26275__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26276__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26277__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26278__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26282__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26283__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26284__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26285__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26286__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26287__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26288__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26289__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26290__RESET_B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__26291__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26293__CLK (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__26293__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26304__RESET_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__26305__RESET_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__26306__RESET_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__26307__RESET_B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__26310__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26311__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26319__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26325__CLK (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__26330__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__26336__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26337__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26340__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26341__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26342__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26343__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26344__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26345__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26346__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26347__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__26350__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26351__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26352__RESET_B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__26362__RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__26529__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26537__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26545__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26553__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26654__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__26657__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__26668__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26670__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26676__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26677__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26684__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26687__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__26692__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26698__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26699__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26700__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26706__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26707__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26708__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26714__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__26743__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26744__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26745__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26746__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26747__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26748__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26749__RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__26750__RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__26861__RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__26862__RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__26875__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__26876__RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__26877__RESET_B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__27053__RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__27065__RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__27067__RESET_B (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__27091__RESET_B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__27093__RESET_B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__27101__RESET_B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__27203__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27210__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27211__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27214__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27218__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27219__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27220__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27221__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27222__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27224__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27226__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27227__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27228__RESET_B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__27230__RESET_B (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__27252__RESET_B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__27259__RESET_B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__27330__RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__27338__RESET_B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__27446__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27451__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27452__RESET_B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__27566__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__27571__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__27574__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__27647__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27648__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27650__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27652__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27653__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27655__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27658__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27661__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27663__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27671__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27680__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27739__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27747__RESET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__27749__RESET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__27750__RESET_B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__27751__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27753__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27755__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27756__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27757__RESET_B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__27762__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27764__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27766__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27767__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27768__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27769__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27770__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27771__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27772__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27773__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27774__RESET_B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__27947__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__27955__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__27990__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__27995__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__27997__RESET_B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__28402__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28407__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28412__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28415__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__28416__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__28417__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28418__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__28420__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28452__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28462__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28466__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28469__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28470__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28471__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28472__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28473__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28474__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28475__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28478__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28482__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__28486__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28487__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28488__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28489__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28491__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28492__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__28495__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28496__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__28497__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28498__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28499__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28504__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28505__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28506__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28507__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28508__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__28513__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28515__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28516__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__28517__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__28519__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__28520__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__28521__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__28602__RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__28721__RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__28729__RESET_B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__28737__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28741__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28742__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28748__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28749__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28750__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28761__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28764__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28765__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28768__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28769__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28770__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28771__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__28796__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28912__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__28919__RESET_B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_0__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_10__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_11__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_12__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_13__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_14__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_15__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_16__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_17__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_18__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_19__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_1__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_20__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_21__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_22__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_23__f_clk_i_A (.DIODE(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_24__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_25__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_26__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_27__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_28__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_29__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_2__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_30__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_31__f_clk_i_A (.DIODE(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_3__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_4__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_5__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_6__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_7__f_clk_i_A (.DIODE(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_8__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_5_9__f_clk_i_A (.DIODE(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_i_A (.DIODE(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_i_A (.DIODE(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_clk_i_A (.DIODE(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_189_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_190_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_191_clk_i_A (.DIODE(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_192_clk_i_A (.DIODE(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_193_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_194_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_195_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_196_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_197_clk_i_A (.DIODE(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_198_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_199_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_200_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_201_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_202_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_203_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_204_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_205_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_206_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_207_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_208_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_209_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_210_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_211_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_212_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_213_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_214_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_215_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_216_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_217_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_218_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_219_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_220_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_221_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_222_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_223_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_224_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_225_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_226_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_227_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_228_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_229_clk_i_A (.DIODE(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_230_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_231_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_232_clk_i_A (.DIODE(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_233_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_234_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_235_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_236_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_237_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_238_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_239_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_240_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_241_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_242_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_243_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_244_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_245_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_246_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_247_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_248_clk_i_A (.DIODE(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_249_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_250_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_251_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_252_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_253_clk_i_A (.DIODE(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_254_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_255_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_256_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_257_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_258_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_259_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_260_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_261_clk_i_A (.DIODE(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_262_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_263_clk_i_A (.DIODE(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_264_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_265_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_266_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_267_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_268_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_269_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_270_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_271_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_272_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_273_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_274_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_275_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_276_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_277_clk_i_A (.DIODE(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_278_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_279_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_280_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_281_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_282_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_283_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_284_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_285_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_286_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_287_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_288_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_289_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_290_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_291_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_292_clk_i_A (.DIODE(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_293_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_294_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_295_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_296_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_297_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_298_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_299_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_300_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_301_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_302_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_303_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_304_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_305_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_306_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_307_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_308_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_309_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_310_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_311_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_312_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_313_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_314_clk_i_A (.DIODE(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_315_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_316_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_317_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_318_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_319_clk_i_A (.DIODE(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_320_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_321_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_322_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_323_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_324_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_325_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_326_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_327_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_328_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_329_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_330_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_331_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_332_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_333_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_334_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_335_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_336_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_337_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_338_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_339_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_340_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_341_clk_i_A (.DIODE(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_342_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_343_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_344_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_345_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_346_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_347_clk_i_A (.DIODE(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_348_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_349_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_350_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_351_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_352_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_353_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_354_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_355_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_356_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_357_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_358_clk_i_A (.DIODE(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_359_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_360_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_361_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_362_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_363_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_364_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_365_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_366_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_367_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_368_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_370_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_371_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_i_A (.DIODE(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_i_A (.DIODE(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_i_A (.DIODE(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_i_A (.DIODE(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_i_A (.DIODE(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_i_A (.DIODE(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_i_A (.DIODE(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_i_A (.DIODE(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_i_A (.DIODE(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_i_A (.DIODE(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_i_A (.DIODE(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_i_A (.DIODE(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_i_A (.DIODE(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3494_A (.DIODE(\line_cache[287][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3508_A (.DIODE(\base_v_bporch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3520_A (.DIODE(\line_cache[287][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3521_A (.DIODE(\res_h_active[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3526_A (.DIODE(\res_h_counter[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3528_A (.DIODE(\line_cache[287][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3530_A (.DIODE(\line_cache[287][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3531_A (.DIODE(\line_cache[287][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3535_A (.DIODE(\line_cache[287][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3536_A (.DIODE(\line_cache[287][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3540_A (.DIODE(\res_h_active[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3541_A (.DIODE(\line_cache[287][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3542_A (.DIODE(\res_h_active[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3575_A (.DIODE(\base_v_bporch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3577_A (.DIODE(\res_h_active[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3578_A (.DIODE(\res_h_active[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3581_A (.DIODE(\res_h_active[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3582_A (.DIODE(\res_h_active[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3585_A (.DIODE(\res_h_active[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3609_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3612_A (.DIODE(\line_cache_idx[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire135_A (.DIODE(_09495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire136_A (.DIODE(_10382_));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _13089_ (.A(net3756),
    .Y(_08829_));
 sky130_fd_sc_hd__nor2_2 _13090_ (.A(\prescaler[0] ),
    .B(net3866),
    .Y(_08830_));
 sky130_fd_sc_hd__inv_2 _13091_ (.A(net3891),
    .Y(_08831_));
 sky130_fd_sc_hd__a311o_1 _13092_ (.A1(_08830_),
    .A2(_08829_),
    .A3(\prescaler_counter[2] ),
    .B1(\prescaler_counter[3] ),
    .C1(_08831_),
    .X(_08832_));
 sky130_fd_sc_hd__or3_1 _13093_ (.A(net3872),
    .B(net4002),
    .C(net3979),
    .X(_08833_));
 sky130_fd_sc_hd__a2111oi_1 _13094_ (.A1(net4000),
    .A2(_08831_),
    .B1(net3984),
    .C1(net3888),
    .D1(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__o311a_1 _13095_ (.A1(\prescaler_counter[2] ),
    .A2(_08829_),
    .A3(_08830_),
    .B1(_08832_),
    .C1(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__inv_2 _13096_ (.A(net4000),
    .Y(_08836_));
 sky130_fd_sc_hd__o21ai_1 _13097_ (.A1(_08829_),
    .A2(_08830_),
    .B1(net3991),
    .Y(_08837_));
 sky130_fd_sc_hd__nand2_1 _13098_ (.A(_08830_),
    .B(_08829_),
    .Y(_08838_));
 sky130_fd_sc_hd__a22o_1 _13099_ (.A1(_08836_),
    .A2(net3891),
    .B1(_08837_),
    .B2(_08838_),
    .X(_08839_));
 sky130_fd_sc_hd__inv_2 _13100_ (.A(net2387),
    .Y(_08840_));
 sky130_fd_sc_hd__nand2_1 _13101_ (.A(_08840_),
    .B(net3952),
    .Y(_08841_));
 sky130_fd_sc_hd__or2_1 _13102_ (.A(net3952),
    .B(_08840_),
    .X(_08842_));
 sky130_fd_sc_hd__nand2_1 _13103_ (.A(\prescaler[0] ),
    .B(\prescaler[1] ),
    .Y(_08843_));
 sky130_fd_sc_hd__or2b_1 _13104_ (.A(_08830_),
    .B_N(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__xor2_1 _13105_ (.A(net3958),
    .B(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__a21o_1 _13106_ (.A1(_08841_),
    .A2(_08842_),
    .B1(_08845_),
    .X(_08846_));
 sky130_fd_sc_hd__inv_2 _13107_ (.A(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__nand3_4 _13108_ (.A(net4003),
    .B(_08839_),
    .C(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nor2_1 _13109_ (.A(\resolution[0] ),
    .B(\resolution[1] ),
    .Y(_08849_));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__nor2_1 _13111_ (.A(\resolution[2] ),
    .B(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__inv_2 _13112_ (.A(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__or2_1 _13113_ (.A(\resolution[3] ),
    .B(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__inv_2 _13114_ (.A(net1999),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(\resolution[0] ),
    .B(\resolution[1] ),
    .Y(_08855_));
 sky130_fd_sc_hd__nand2_1 _13116_ (.A(_08850_),
    .B(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__or2_1 _13117_ (.A(_08854_),
    .B(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__nand2_1 _13118_ (.A(_08856_),
    .B(_08854_),
    .Y(_08858_));
 sky130_fd_sc_hd__xor2_1 _13119_ (.A(\pixel_double_counter[0] ),
    .B(\resolution[0] ),
    .X(_08859_));
 sky130_fd_sc_hd__and4_1 _13120_ (.A(_08853_),
    .B(_08857_),
    .C(_08858_),
    .D(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__inv_2 _13121_ (.A(net1862),
    .Y(_08861_));
 sky130_fd_sc_hd__nand2_1 _13122_ (.A(_08852_),
    .B(net3738),
    .Y(_08862_));
 sky130_fd_sc_hd__nand2_1 _13123_ (.A(_08853_),
    .B(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__xor2_1 _13124_ (.A(_08861_),
    .B(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__inv_2 _13125_ (.A(net1940),
    .Y(_08865_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(_08850_),
    .B(\resolution[2] ),
    .Y(_08866_));
 sky130_fd_sc_hd__nand2_1 _13127_ (.A(_08852_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__xor2_1 _13128_ (.A(_08865_),
    .B(_08867_),
    .X(_08868_));
 sky130_fd_sc_hd__and3_1 _13129_ (.A(_08860_),
    .B(_08864_),
    .C(_08868_),
    .X(_08869_));
 sky130_fd_sc_hd__inv_2 _13130_ (.A(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__inv_2 _13131_ (.A(net3990),
    .Y(_08871_));
 sky130_fd_sc_hd__inv_2 _13132_ (.A(\base_h_active[7] ),
    .Y(_08872_));
 sky130_fd_sc_hd__nor2_1 _13133_ (.A(\base_h_counter[7] ),
    .B(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__inv_2 _13134_ (.A(net3968),
    .Y(_08874_));
 sky130_fd_sc_hd__nor2_1 _13135_ (.A(\base_h_active[7] ),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__inv_2 _13136_ (.A(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__o21ai_1 _13137_ (.A1(_08871_),
    .A2(\base_h_active[6] ),
    .B1(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__a211oi_1 _13138_ (.A1(_08871_),
    .A2(\base_h_active[6] ),
    .B1(_08873_),
    .C1(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__inv_2 _13139_ (.A(net3994),
    .Y(_08879_));
 sky130_fd_sc_hd__nand2_1 _13140_ (.A(_08879_),
    .B(\base_h_active[4] ),
    .Y(_08880_));
 sky130_fd_sc_hd__inv_2 _13141_ (.A(\base_h_active[4] ),
    .Y(_08881_));
 sky130_fd_sc_hd__nand2_1 _13142_ (.A(_08881_),
    .B(\base_h_counter[4] ),
    .Y(_08882_));
 sky130_fd_sc_hd__inv_2 _13143_ (.A(\base_h_active[5] ),
    .Y(_08883_));
 sky130_fd_sc_hd__nor2_1 _13144_ (.A(\base_h_counter[5] ),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__inv_2 _13145_ (.A(net3992),
    .Y(_08885_));
 sky130_fd_sc_hd__nor2_1 _13146_ (.A(\base_h_active[5] ),
    .B(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__nor2_1 _13147_ (.A(_08884_),
    .B(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__and4_2 _13148_ (.A(_08878_),
    .B(_08880_),
    .C(_08882_),
    .D(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__inv_2 _13149_ (.A(\base_h_active[0] ),
    .Y(_08889_));
 sky130_fd_sc_hd__inv_2 _13150_ (.A(net1985),
    .Y(_08890_));
 sky130_fd_sc_hd__inv_2 _13151_ (.A(net3965),
    .Y(_08891_));
 sky130_fd_sc_hd__nand2_1 _13152_ (.A(_08891_),
    .B(\base_h_active[1] ),
    .Y(_08892_));
 sky130_fd_sc_hd__inv_2 _13153_ (.A(\base_h_active[1] ),
    .Y(_08893_));
 sky130_fd_sc_hd__nand2_1 _13154_ (.A(_08893_),
    .B(\base_h_counter[1] ),
    .Y(_08894_));
 sky130_fd_sc_hd__o211a_1 _13155_ (.A1(\base_h_active[0] ),
    .A2(_08890_),
    .B1(_08892_),
    .C1(_08894_),
    .X(_08895_));
 sky130_fd_sc_hd__inv_2 _13156_ (.A(\base_h_active[2] ),
    .Y(_08896_));
 sky130_fd_sc_hd__nor2_1 _13157_ (.A(\base_h_counter[2] ),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__inv_2 _13158_ (.A(net3976),
    .Y(_08898_));
 sky130_fd_sc_hd__nor2_1 _13159_ (.A(\base_h_active[2] ),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__nor2_1 _13160_ (.A(_08897_),
    .B(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__inv_2 _13161_ (.A(net3988),
    .Y(_08901_));
 sky130_fd_sc_hd__nand2_1 _13162_ (.A(_08901_),
    .B(\base_h_active[3] ),
    .Y(_08902_));
 sky130_fd_sc_hd__inv_2 _13163_ (.A(\base_h_active[3] ),
    .Y(_08903_));
 sky130_fd_sc_hd__nand2_1 _13164_ (.A(_08903_),
    .B(\base_h_counter[3] ),
    .Y(_08904_));
 sky130_fd_sc_hd__and3_1 _13165_ (.A(_08900_),
    .B(_08902_),
    .C(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__inv_2 _13166_ (.A(\base_h_active[9] ),
    .Y(_08906_));
 sky130_fd_sc_hd__nor2_1 _13167_ (.A(net3947),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(_08906_),
    .B(\base_h_counter[9] ),
    .Y(_08908_));
 sky130_fd_sc_hd__and2b_1 _13169_ (.A_N(_08907_),
    .B(_08908_),
    .X(_08909_));
 sky130_fd_sc_hd__inv_2 _13170_ (.A(net3959),
    .Y(_08910_));
 sky130_fd_sc_hd__nand2_1 _13171_ (.A(_08910_),
    .B(\base_h_active[8] ),
    .Y(_08911_));
 sky130_fd_sc_hd__or2_1 _13172_ (.A(\base_h_active[8] ),
    .B(_08910_),
    .X(_08912_));
 sky130_fd_sc_hd__and3_1 _13173_ (.A(_08909_),
    .B(_08911_),
    .C(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__o2111a_1 _13174_ (.A1(_08889_),
    .A2(\base_h_counter[0] ),
    .B1(_08895_),
    .C1(_08905_),
    .D1(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__inv_2 _13175_ (.A(\base_v_active[6] ),
    .Y(_08915_));
 sky130_fd_sc_hd__nor2_1 _13176_ (.A(\base_v_counter[6] ),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__inv_2 _13177_ (.A(\base_v_counter[6] ),
    .Y(_08917_));
 sky130_fd_sc_hd__nor2_1 _13178_ (.A(\base_v_active[6] ),
    .B(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__buf_2 _13179_ (.A(net3936),
    .X(_08919_));
 sky130_fd_sc_hd__inv_2 _13180_ (.A(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__nand2_1 _13181_ (.A(_08920_),
    .B(\base_v_active[7] ),
    .Y(_08921_));
 sky130_fd_sc_hd__inv_2 _13182_ (.A(\base_v_active[7] ),
    .Y(_08922_));
 sky130_fd_sc_hd__nand2_1 _13183_ (.A(_08922_),
    .B(_08919_),
    .Y(_08923_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(_08921_),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__or3_1 _13185_ (.A(_08916_),
    .B(_08918_),
    .C(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__inv_2 _13186_ (.A(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__inv_2 _13187_ (.A(\base_v_active[5] ),
    .Y(_08927_));
 sky130_fd_sc_hd__nor2_1 _13188_ (.A(\base_v_counter[5] ),
    .B(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__inv_2 _13189_ (.A(net3817),
    .Y(_08929_));
 sky130_fd_sc_hd__nor2_1 _13190_ (.A(\base_v_active[5] ),
    .B(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__nor2_1 _13191_ (.A(_08928_),
    .B(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__inv_2 _13192_ (.A(\base_v_active[4] ),
    .Y(_08932_));
 sky130_fd_sc_hd__nor2_1 _13193_ (.A(\base_v_counter[4] ),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__inv_2 _13194_ (.A(net3797),
    .Y(_08934_));
 sky130_fd_sc_hd__nor2_1 _13195_ (.A(\base_v_active[4] ),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__nor2_1 _13196_ (.A(_08933_),
    .B(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__and3_2 _13197_ (.A(_08926_),
    .B(_08931_),
    .C(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__inv_2 _13198_ (.A(net2025),
    .Y(_08938_));
 sky130_fd_sc_hd__inv_2 _13199_ (.A(\base_v_active[8] ),
    .Y(_08939_));
 sky130_fd_sc_hd__nor2_1 _13200_ (.A(\base_v_counter[8] ),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__inv_2 _13201_ (.A(\base_v_counter[8] ),
    .Y(_08941_));
 sky130_fd_sc_hd__nor2_1 _13202_ (.A(\base_v_active[8] ),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__or3_2 _13203_ (.A(\base_v_counter[9] ),
    .B(_08940_),
    .C(_08942_),
    .X(_08943_));
 sky130_fd_sc_hd__inv_2 _13204_ (.A(net3784),
    .Y(_08944_));
 sky130_fd_sc_hd__nand2_1 _13205_ (.A(_08944_),
    .B(\base_v_active[3] ),
    .Y(_08945_));
 sky130_fd_sc_hd__inv_2 _13206_ (.A(\base_v_active[3] ),
    .Y(_08946_));
 sky130_fd_sc_hd__nand2_1 _13207_ (.A(_08946_),
    .B(\base_v_counter[3] ),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_1 _13208_ (.A(_08945_),
    .B(_08947_),
    .Y(_08948_));
 sky130_fd_sc_hd__inv_2 _13209_ (.A(net2011),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_1 _13210_ (.A(_08949_),
    .B(\base_v_active[2] ),
    .Y(_08950_));
 sky130_fd_sc_hd__or2_1 _13211_ (.A(\base_v_active[2] ),
    .B(_08949_),
    .X(_08951_));
 sky130_fd_sc_hd__and3b_1 _13212_ (.A_N(_08948_),
    .B(_08950_),
    .C(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__inv_2 _13213_ (.A(\base_v_active[1] ),
    .Y(_08953_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(\base_v_counter[1] ),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_1 _13215_ (.A(_08953_),
    .B(\base_v_counter[1] ),
    .Y(_08955_));
 sky130_fd_sc_hd__o21ai_1 _13216_ (.A1(\base_v_active[0] ),
    .A2(_08938_),
    .B1(_08955_),
    .Y(_08956_));
 sky130_fd_sc_hd__nor2_1 _13217_ (.A(_08954_),
    .B(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__nand2_1 _13218_ (.A(_08952_),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__a211oi_4 _13219_ (.A1(\base_v_active[0] ),
    .A2(_08938_),
    .B1(_08943_),
    .C1(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__inv_2 _13220_ (.A(net3713),
    .Y(_08960_));
 sky130_fd_sc_hd__a21o_1 _13221_ (.A1(_08931_),
    .A2(_08933_),
    .B1(_08928_),
    .X(_08961_));
 sky130_fd_sc_hd__or2_1 _13222_ (.A(_08954_),
    .B(_08957_),
    .X(_08962_));
 sky130_fd_sc_hd__o21ai_1 _13223_ (.A1(_08950_),
    .A2(_08948_),
    .B1(_08945_),
    .Y(_08963_));
 sky130_fd_sc_hd__a21o_1 _13224_ (.A1(_08952_),
    .A2(_08962_),
    .B1(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__a21bo_1 _13225_ (.A1(_08923_),
    .A2(_08916_),
    .B1_N(_08921_),
    .X(_08965_));
 sky130_fd_sc_hd__a221oi_2 _13226_ (.A1(_08926_),
    .A2(_08961_),
    .B1(_08937_),
    .B2(_08964_),
    .C1(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__o2bb2a_1 _13227_ (.A1_N(_08960_),
    .A2_N(_08940_),
    .B1(_08943_),
    .B2(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__a221oi_4 _13228_ (.A1(_08888_),
    .A2(_08914_),
    .B1(_08937_),
    .B2(_08959_),
    .C1(_08967_),
    .Y(_08968_));
 sky130_fd_sc_hd__a31o_1 _13229_ (.A1(_08887_),
    .A2(\base_h_active[4] ),
    .A3(_08879_),
    .B1(_08884_),
    .X(_08969_));
 sky130_fd_sc_hd__or2b_1 _13230_ (.A(_08895_),
    .B_N(_08892_),
    .X(_08970_));
 sky130_fd_sc_hd__and3_1 _13231_ (.A(_08897_),
    .B(_08902_),
    .C(_08904_),
    .X(_08971_));
 sky130_fd_sc_hd__a221o_1 _13232_ (.A1(_08901_),
    .A2(\base_h_active[3] ),
    .B1(_08970_),
    .B2(_08905_),
    .C1(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__a31o_1 _13233_ (.A1(_08876_),
    .A2(_08871_),
    .A3(\base_h_active[6] ),
    .B1(_08873_),
    .X(_08973_));
 sky130_fd_sc_hd__a221o_1 _13234_ (.A1(_08878_),
    .A2(_08969_),
    .B1(_08972_),
    .B2(_08888_),
    .C1(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__a31o_1 _13235_ (.A1(_08908_),
    .A2(_08910_),
    .A3(\base_h_active[8] ),
    .B1(_08907_),
    .X(_08975_));
 sky130_fd_sc_hd__a21o_1 _13236_ (.A1(_08974_),
    .A2(_08913_),
    .B1(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__nand2_2 _13237_ (.A(_08968_),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__inv_2 _13238_ (.A(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__nand2_8 _13239_ (.A(_08978_),
    .B(net49),
    .Y(_08979_));
 sky130_fd_sc_hd__nor3_1 _13240_ (.A(_08848_),
    .B(_08870_),
    .C(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__inv_2 _13241_ (.A(net2797),
    .Y(_08981_));
 sky130_fd_sc_hd__nand2_1 _13242_ (.A(_08856_),
    .B(_08981_),
    .Y(_08982_));
 sky130_fd_sc_hd__or2_1 _13243_ (.A(_08981_),
    .B(_08856_),
    .X(_08983_));
 sky130_fd_sc_hd__xor2_1 _13244_ (.A(\resolution[0] ),
    .B(\line_double_counter[0] ),
    .X(_08984_));
 sky130_fd_sc_hd__and4_1 _13245_ (.A(_08853_),
    .B(_08982_),
    .C(_08983_),
    .D(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__inv_2 _13246_ (.A(net1992),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_1 _13247_ (.A(_08867_),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__or2_1 _13248_ (.A(_08986_),
    .B(_08867_),
    .X(_08988_));
 sky130_fd_sc_hd__and3_1 _13249_ (.A(_08985_),
    .B(_08987_),
    .C(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__xor2_1 _13250_ (.A(net2005),
    .B(_08863_),
    .X(_08990_));
 sky130_fd_sc_hd__inv_2 _13251_ (.A(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__nand2_1 _13252_ (.A(_08989_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__clkbuf_16 _13253_ (.A(\res_h_counter[8] ),
    .X(_08993_));
 sky130_fd_sc_hd__inv_4 _13254_ (.A(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__clkbuf_16 _13255_ (.A(_08994_),
    .X(_08995_));
 sky130_fd_sc_hd__nor2_1 _13256_ (.A(\res_h_active[8] ),
    .B(_08995_),
    .Y(_08996_));
 sky130_fd_sc_hd__and2_1 _13257_ (.A(_08995_),
    .B(\res_h_active[8] ),
    .X(_08997_));
 sky130_fd_sc_hd__nor2_1 _13258_ (.A(_08996_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__nor2_1 _13259_ (.A(\res_h_active[2] ),
    .B(\res_h_active[3] ),
    .Y(_08999_));
 sky130_fd_sc_hd__clkinvlp_2 _13260_ (.A(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__nor2_1 _13261_ (.A(\res_h_active[0] ),
    .B(\res_h_active[1] ),
    .Y(_09001_));
 sky130_fd_sc_hd__inv_2 _13262_ (.A(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__nor2_1 _13263_ (.A(_09000_),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__inv_2 _13264_ (.A(\res_h_active[4] ),
    .Y(_09004_));
 sky130_fd_sc_hd__nand2_1 _13265_ (.A(_09003_),
    .B(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__or2_1 _13266_ (.A(\res_h_active[5] ),
    .B(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__nor2_1 _13267_ (.A(\res_h_active[6] ),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__inv_2 _13268_ (.A(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__nor2_1 _13269_ (.A(\res_h_active[7] ),
    .B(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(_08998_),
    .A1(_08997_),
    .S(_09009_),
    .X(_09010_));
 sky130_fd_sc_hd__nand2_1 _13271_ (.A(_09006_),
    .B(net3970),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_1 _13272_ (.A(_09008_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__inv_6 _13273_ (.A(net1997),
    .Y(_09013_));
 sky130_fd_sc_hd__nand2_1 _13274_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__xnor2_1 _13275_ (.A(\res_h_active[1] ),
    .B(\res_h_counter[1] ),
    .Y(_09015_));
 sky130_fd_sc_hd__inv_2 _13276_ (.A(net1959),
    .Y(_09016_));
 sky130_fd_sc_hd__inv_2 _13277_ (.A(net3773),
    .Y(_09017_));
 sky130_fd_sc_hd__nand2_1 _13278_ (.A(_09017_),
    .B(\res_h_active[0] ),
    .Y(_09018_));
 sky130_fd_sc_hd__o21ai_1 _13279_ (.A1(\res_h_active[0] ),
    .A2(_09015_),
    .B1(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__o211a_1 _13280_ (.A1(\res_h_counter[0] ),
    .A2(_09015_),
    .B1(_09016_),
    .C1(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__inv_2 _13281_ (.A(net3638),
    .Y(_09021_));
 sky130_fd_sc_hd__or2_1 _13282_ (.A(\res_h_active[2] ),
    .B(_09002_),
    .X(_09022_));
 sky130_fd_sc_hd__nand2_1 _13283_ (.A(_09022_),
    .B(\res_h_active[3] ),
    .Y(_09023_));
 sky130_fd_sc_hd__inv_2 _13284_ (.A(_09003_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__or2_1 _13286_ (.A(_09021_),
    .B(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__nand2_1 _13287_ (.A(_09002_),
    .B(\res_h_active[2] ),
    .Y(_09027_));
 sky130_fd_sc_hd__nand2_1 _13288_ (.A(_09022_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__inv_2 _13289_ (.A(net3745),
    .Y(_09029_));
 sky130_fd_sc_hd__nand2_1 _13290_ (.A(_09028_),
    .B(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__or2_1 _13291_ (.A(_09029_),
    .B(_09028_),
    .X(_09031_));
 sky130_fd_sc_hd__nand2_1 _13292_ (.A(_09025_),
    .B(_09021_),
    .Y(_09032_));
 sky130_fd_sc_hd__and4_1 _13293_ (.A(_09026_),
    .B(_09030_),
    .C(_09031_),
    .D(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__and4_1 _13294_ (.A(_09010_),
    .B(_09014_),
    .C(_09020_),
    .D(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__inv_2 _13295_ (.A(net3915),
    .Y(_09035_));
 sky130_fd_sc_hd__and2_1 _13296_ (.A(_09008_),
    .B(\res_h_active[7] ),
    .X(_09036_));
 sky130_fd_sc_hd__or2_1 _13297_ (.A(_09009_),
    .B(_09036_),
    .X(_09037_));
 sky130_fd_sc_hd__or2_1 _13298_ (.A(_09035_),
    .B(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__nand2_1 _13299_ (.A(_09037_),
    .B(_09035_),
    .Y(_09039_));
 sky130_fd_sc_hd__and3_2 _13300_ (.A(_09034_),
    .B(_09038_),
    .C(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__nand2_1 _13301_ (.A(_09005_),
    .B(\res_h_active[5] ),
    .Y(_09041_));
 sky130_fd_sc_hd__nand2_1 _13302_ (.A(_09006_),
    .B(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__inv_2 _13303_ (.A(net3902),
    .Y(_09043_));
 sky130_fd_sc_hd__nand2_1 _13304_ (.A(_09042_),
    .B(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__nand2_1 _13305_ (.A(_09024_),
    .B(\res_h_active[4] ),
    .Y(_09045_));
 sky130_fd_sc_hd__nand2_1 _13306_ (.A(_09045_),
    .B(_09005_),
    .Y(_09046_));
 sky130_fd_sc_hd__inv_2 _13307_ (.A(net3943),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_1 _13308_ (.A(_09046_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__or2_1 _13309_ (.A(_09047_),
    .B(_09046_),
    .X(_09049_));
 sky130_fd_sc_hd__o211a_1 _13310_ (.A1(_09043_),
    .A2(_09042_),
    .B1(_09048_),
    .C1(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__o211a_1 _13311_ (.A1(_09013_),
    .A2(_09012_),
    .B1(_09044_),
    .C1(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__nand2_8 _13312_ (.A(_09040_),
    .B(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__or2_1 _13313_ (.A(_08992_),
    .B(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__nand2_1 _13314_ (.A(_08980_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__nor2_1 _13315_ (.A(_08848_),
    .B(_08977_),
    .Y(_09055_));
 sky130_fd_sc_hd__inv_2 _13316_ (.A(net49),
    .Y(_09056_));
 sky130_fd_sc_hd__buf_12 _13317_ (.A(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__a21o_1 _13318_ (.A1(_09055_),
    .A2(_08869_),
    .B1(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__inv_2 _13319_ (.A(net1994),
    .Y(_09059_));
 sky130_fd_sc_hd__a21o_1 _13320_ (.A1(_09054_),
    .A2(_09058_),
    .B1(_09059_),
    .X(_09060_));
 sky130_fd_sc_hd__nand2_1 _13321_ (.A(_08999_),
    .B(_09004_),
    .Y(_09061_));
 sky130_fd_sc_hd__nor2_1 _13322_ (.A(\res_h_active[5] ),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__inv_2 _13323_ (.A(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nor2_1 _13324_ (.A(\res_h_active[6] ),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__inv_2 _13325_ (.A(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__nor2_1 _13326_ (.A(net3966),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__inv_2 _13327_ (.A(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(_09065_),
    .B(net3966),
    .Y(_09068_));
 sky130_fd_sc_hd__and2_1 _13329_ (.A(_09067_),
    .B(_09068_),
    .X(_09069_));
 sky130_fd_sc_hd__buf_8 _13330_ (.A(\line_cache_idx[8] ),
    .X(_09070_));
 sky130_fd_sc_hd__inv_2 _13331_ (.A(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__nor2_1 _13332_ (.A(net3971),
    .B(_09067_),
    .Y(_09072_));
 sky130_fd_sc_hd__inv_2 _13333_ (.A(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__nand2_1 _13334_ (.A(_09067_),
    .B(net3971),
    .Y(_09074_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(_09073_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__or2_1 _13336_ (.A(_09071_),
    .B(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__inv_2 _13337_ (.A(net3989),
    .Y(_09077_));
 sky130_fd_sc_hd__nand2_1 _13338_ (.A(_09075_),
    .B(_09071_),
    .Y(_09078_));
 sky130_fd_sc_hd__and4_1 _13339_ (.A(_09076_),
    .B(_09077_),
    .C(_09073_),
    .D(_09078_),
    .X(_09079_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_09063_),
    .B(\res_h_active[6] ),
    .Y(_09080_));
 sky130_fd_sc_hd__inv_2 _13341_ (.A(net3921),
    .Y(_09081_));
 sky130_fd_sc_hd__nand2_1 _13342_ (.A(\res_h_active[2] ),
    .B(\res_h_active[3] ),
    .Y(_09082_));
 sky130_fd_sc_hd__nand2_1 _13343_ (.A(_09000_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__o21ai_1 _13344_ (.A1(\line_cache_idx[2] ),
    .A2(_09001_),
    .B1(\res_h_active[2] ),
    .Y(_09084_));
 sky130_fd_sc_hd__nand2_1 _13345_ (.A(_09001_),
    .B(\line_cache_idx[2] ),
    .Y(_09085_));
 sky130_fd_sc_hd__a22o_1 _13346_ (.A1(_09083_),
    .A2(_09081_),
    .B1(_09084_),
    .B2(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__o21ai_1 _13347_ (.A1(_09081_),
    .A2(_09083_),
    .B1(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__nand2_1 _13348_ (.A(_09000_),
    .B(\res_h_active[4] ),
    .Y(_09088_));
 sky130_fd_sc_hd__nand2_1 _13349_ (.A(_09088_),
    .B(_09061_),
    .Y(_09089_));
 sky130_fd_sc_hd__inv_2 _13350_ (.A(net3995),
    .Y(_09090_));
 sky130_fd_sc_hd__nand2_1 _13351_ (.A(_09089_),
    .B(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__inv_2 _13352_ (.A(net3381),
    .Y(_09092_));
 sky130_fd_sc_hd__nand2_1 _13353_ (.A(_09061_),
    .B(\res_h_active[5] ),
    .Y(_09093_));
 sky130_fd_sc_hd__nand2_1 _13354_ (.A(_09063_),
    .B(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__o22ai_1 _13355_ (.A1(_09090_),
    .A2(_09089_),
    .B1(_09092_),
    .B2(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__a21o_1 _13356_ (.A1(_09087_),
    .A2(_09091_),
    .B1(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__a21o_1 _13357_ (.A1(_09065_),
    .A2(_09080_),
    .B1(\line_cache_idx[6] ),
    .X(_09097_));
 sky130_fd_sc_hd__nand2_1 _13358_ (.A(_09094_),
    .B(_09092_),
    .Y(_09098_));
 sky130_fd_sc_hd__and3_1 _13359_ (.A(_09096_),
    .B(_09097_),
    .C(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__a31o_1 _13360_ (.A1(\line_cache_idx[6] ),
    .A2(_09065_),
    .A3(_09080_),
    .B1(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__a31o_1 _13361_ (.A1(net3913),
    .A2(_09067_),
    .A3(_09068_),
    .B1(_09100_),
    .X(_09101_));
 sky130_fd_sc_hd__o211ai_2 _13362_ (.A1(net3913),
    .A2(_09069_),
    .B1(_09079_),
    .C1(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__and4_1 _13363_ (.A(_09073_),
    .B(_09074_),
    .C(_09070_),
    .D(_09077_),
    .X(_09103_));
 sky130_fd_sc_hd__a21oi_1 _13364_ (.A1(net3989),
    .A2(_09073_),
    .B1(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__nand2_4 _13365_ (.A(_09102_),
    .B(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__buf_6 _13366_ (.A(net3972),
    .X(_09106_));
 sky130_fd_sc_hd__inv_4 _13367_ (.A(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__nand2_2 _13368_ (.A(net49),
    .B(net75),
    .Y(_09108_));
 sky130_fd_sc_hd__nor2_8 _13369_ (.A(_09107_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__clkbuf_16 _13370_ (.A(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__nand2_4 _13371_ (.A(_09105_),
    .B(_09110_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand2_1 _13372_ (.A(net1995),
    .B(_09111_),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _13373_ (.A(_09105_),
    .Y(_09112_));
 sky130_fd_sc_hd__inv_2 _13374_ (.A(_09108_),
    .Y(_09113_));
 sky130_fd_sc_hd__inv_2 _13375_ (.A(_08848_),
    .Y(_09114_));
 sky130_fd_sc_hd__nor2_1 _13376_ (.A(net75),
    .B(_09057_),
    .Y(_09115_));
 sky130_fd_sc_hd__a31o_1 _13377_ (.A1(_09112_),
    .A2(_09113_),
    .A3(_09114_),
    .B1(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__or2_1 _13378_ (.A(_08992_),
    .B(_08848_),
    .X(_09117_));
 sky130_fd_sc_hd__nor2_1 _13379_ (.A(_08870_),
    .B(_09052_),
    .Y(_09118_));
 sky130_fd_sc_hd__nand2_1 _13380_ (.A(_08978_),
    .B(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__a21o_1 _13381_ (.A1(_09115_),
    .A2(_09117_),
    .B1(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__and3_1 _13382_ (.A(_09116_),
    .B(_09120_),
    .C(_09106_),
    .X(_09121_));
 sky130_fd_sc_hd__and3_1 _13383_ (.A(_09118_),
    .B(_09106_),
    .C(_08992_),
    .X(_09122_));
 sky130_fd_sc_hd__a32o_1 _13384_ (.A1(_09055_),
    .A2(_09122_),
    .A3(_09113_),
    .B1(_09110_),
    .B2(_08848_),
    .X(_09123_));
 sky130_fd_sc_hd__nand2_1 _13385_ (.A(_09123_),
    .B(_09112_),
    .Y(_09124_));
 sky130_fd_sc_hd__clkbuf_16 _13386_ (.A(net49),
    .X(_09125_));
 sky130_fd_sc_hd__clkbuf_16 _13387_ (.A(_09125_),
    .X(_09126_));
 sky130_fd_sc_hd__buf_8 _13388_ (.A(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__nand2_4 _13389_ (.A(_09127_),
    .B(net3977),
    .Y(_09128_));
 sky130_fd_sc_hd__nand3b_1 _13390_ (.A_N(_09121_),
    .B(_09124_),
    .C(_09128_),
    .Y(_00010_));
 sky130_fd_sc_hd__buf_8 _13391_ (.A(_09057_),
    .X(_09129_));
 sky130_fd_sc_hd__buf_8 _13392_ (.A(_09129_),
    .X(_09130_));
 sky130_fd_sc_hd__inv_2 _13393_ (.A(_09055_),
    .Y(_09131_));
 sky130_fd_sc_hd__a211oi_1 _13394_ (.A1(net75),
    .A2(_09105_),
    .B1(_09130_),
    .C1(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__nor2_2 _13395_ (.A(_08870_),
    .B(_09053_),
    .Y(_09133_));
 sky130_fd_sc_hd__nor2_1 _13396_ (.A(_09059_),
    .B(_09053_),
    .Y(_09134_));
 sky130_fd_sc_hd__a21o_1 _13397_ (.A1(_08980_),
    .A2(_09134_),
    .B1(_09130_),
    .X(_09135_));
 sky130_fd_sc_hd__a31o_1 _13398_ (.A1(_09106_),
    .A2(_09132_),
    .A3(_09133_),
    .B1(_09135_),
    .X(_00011_));
 sky130_fd_sc_hd__inv_2 _13399_ (.A(\base_h_fporch[3] ),
    .Y(_09136_));
 sky130_fd_sc_hd__nand2_1 _13400_ (.A(_08903_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__nand2_1 _13401_ (.A(\base_h_active[3] ),
    .B(\base_h_fporch[3] ),
    .Y(_09138_));
 sky130_fd_sc_hd__nand2_1 _13402_ (.A(_09137_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__inv_2 _13403_ (.A(\base_h_fporch[2] ),
    .Y(_09140_));
 sky130_fd_sc_hd__nand2_1 _13404_ (.A(_08896_),
    .B(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__nand2_1 _13405_ (.A(\base_h_active[2] ),
    .B(\base_h_fporch[2] ),
    .Y(_09142_));
 sky130_fd_sc_hd__nand2_1 _13406_ (.A(_09141_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__nor2_1 _13407_ (.A(_09139_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__nand2_1 _13408_ (.A(\base_h_active[0] ),
    .B(\base_h_fporch[0] ),
    .Y(_09145_));
 sky130_fd_sc_hd__nor2_1 _13409_ (.A(\base_h_active[1] ),
    .B(\base_h_fporch[1] ),
    .Y(_09146_));
 sky130_fd_sc_hd__nand2_1 _13410_ (.A(\base_h_active[1] ),
    .B(\base_h_fporch[1] ),
    .Y(_09147_));
 sky130_fd_sc_hd__o21ai_1 _13411_ (.A1(_09145_),
    .A2(_09146_),
    .B1(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__nand2_1 _13412_ (.A(_09144_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__nor2_1 _13413_ (.A(\base_h_active[3] ),
    .B(\base_h_fporch[3] ),
    .Y(_09150_));
 sky130_fd_sc_hd__o21a_1 _13414_ (.A1(_09142_),
    .A2(_09150_),
    .B1(_09138_),
    .X(_09151_));
 sky130_fd_sc_hd__nand2_1 _13415_ (.A(_09149_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__or2_1 _13416_ (.A(\base_h_active[4] ),
    .B(\base_h_fporch[4] ),
    .X(_09153_));
 sky130_fd_sc_hd__nand2_1 _13417_ (.A(\base_h_active[4] ),
    .B(\base_h_fporch[4] ),
    .Y(_09154_));
 sky130_fd_sc_hd__nand2_1 _13418_ (.A(_09153_),
    .B(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__inv_2 _13419_ (.A(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__nand2_1 _13420_ (.A(_09156_),
    .B(\base_h_active[5] ),
    .Y(_09157_));
 sky130_fd_sc_hd__inv_2 _13421_ (.A(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(_09152_),
    .B(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__nor2_1 _13423_ (.A(_08883_),
    .B(_09154_),
    .Y(_09160_));
 sky130_fd_sc_hd__inv_2 _13424_ (.A(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__nand2_1 _13425_ (.A(_09159_),
    .B(_09161_),
    .Y(_09162_));
 sky130_fd_sc_hd__nand2_1 _13426_ (.A(_09162_),
    .B(\base_h_active[6] ),
    .Y(_09163_));
 sky130_fd_sc_hd__or2_1 _13427_ (.A(_08872_),
    .B(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__inv_2 _13428_ (.A(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__or2_1 _13429_ (.A(\base_h_active[8] ),
    .B(_09165_),
    .X(_09166_));
 sky130_fd_sc_hd__nand2_1 _13430_ (.A(_09165_),
    .B(\base_h_active[8] ),
    .Y(_09167_));
 sky130_fd_sc_hd__nand2_1 _13431_ (.A(_09166_),
    .B(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__nand2_1 _13432_ (.A(_09163_),
    .B(_08872_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand2_1 _13433_ (.A(_09164_),
    .B(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__a21oi_2 _13434_ (.A1(_09152_),
    .A2(_09158_),
    .B1(_09160_),
    .Y(_09171_));
 sky130_fd_sc_hd__inv_2 _13435_ (.A(\base_h_active[6] ),
    .Y(_09172_));
 sky130_fd_sc_hd__nand2_1 _13436_ (.A(_09171_),
    .B(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__nand2_1 _13437_ (.A(_09173_),
    .B(_09163_),
    .Y(_09174_));
 sky130_fd_sc_hd__inv_2 _13438_ (.A(\base_h_sync[6] ),
    .Y(_09175_));
 sky130_fd_sc_hd__nand2_1 _13439_ (.A(_09174_),
    .B(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__nand3_1 _13440_ (.A(_09173_),
    .B(\base_h_sync[6] ),
    .C(_09163_),
    .Y(_09177_));
 sky130_fd_sc_hd__nand2_1 _13441_ (.A(_09176_),
    .B(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__nor2_1 _13442_ (.A(_09170_),
    .B(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_1 _13443_ (.A(_09152_),
    .B(_09156_),
    .Y(_09180_));
 sky130_fd_sc_hd__nand3_1 _13444_ (.A(_09180_),
    .B(_08883_),
    .C(_09154_),
    .Y(_09181_));
 sky130_fd_sc_hd__nand2_2 _13445_ (.A(_09181_),
    .B(_09171_),
    .Y(_09182_));
 sky130_fd_sc_hd__inv_2 _13446_ (.A(\base_h_sync[5] ),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_1 _13447_ (.A(_09182_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__nand3_1 _13448_ (.A(_09149_),
    .B(_09151_),
    .C(_09155_),
    .Y(_09185_));
 sky130_fd_sc_hd__nand2_1 _13449_ (.A(_09180_),
    .B(_09185_),
    .Y(_09186_));
 sky130_fd_sc_hd__inv_2 _13450_ (.A(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__nand2_1 _13451_ (.A(_09187_),
    .B(\base_h_sync[4] ),
    .Y(_09188_));
 sky130_fd_sc_hd__inv_2 _13452_ (.A(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__nor2_1 _13453_ (.A(_09183_),
    .B(_09182_),
    .Y(_09190_));
 sky130_fd_sc_hd__a21oi_2 _13454_ (.A1(_09184_),
    .A2(_09189_),
    .B1(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__inv_2 _13455_ (.A(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__nand2_1 _13456_ (.A(_09179_),
    .B(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__or2_1 _13457_ (.A(_09177_),
    .B(_09170_),
    .X(_09194_));
 sky130_fd_sc_hd__nand2_1 _13458_ (.A(_09193_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__inv_2 _13459_ (.A(_09145_),
    .Y(_09196_));
 sky130_fd_sc_hd__inv_2 _13460_ (.A(\base_h_fporch[1] ),
    .Y(_09197_));
 sky130_fd_sc_hd__nand2_1 _13461_ (.A(_08893_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand3_2 _13462_ (.A(_09196_),
    .B(_09198_),
    .C(_09147_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand2_1 _13463_ (.A(_08893_),
    .B(\base_h_fporch[1] ),
    .Y(_09200_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(_09197_),
    .B(\base_h_active[1] ),
    .Y(_09201_));
 sky130_fd_sc_hd__nand3_1 _13465_ (.A(_09200_),
    .B(_09201_),
    .C(_09145_),
    .Y(_09202_));
 sky130_fd_sc_hd__nand2_1 _13466_ (.A(_09199_),
    .B(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__inv_2 _13467_ (.A(\base_h_sync[1] ),
    .Y(_09204_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(_09203_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__nand3_1 _13469_ (.A(_09199_),
    .B(_09202_),
    .C(\base_h_sync[1] ),
    .Y(_09206_));
 sky130_fd_sc_hd__nor2_1 _13470_ (.A(\base_h_active[0] ),
    .B(\base_h_fporch[0] ),
    .Y(_09207_));
 sky130_fd_sc_hd__nor2_1 _13471_ (.A(_09207_),
    .B(_09196_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand2_1 _13472_ (.A(_09208_),
    .B(\base_h_sync[0] ),
    .Y(_09209_));
 sky130_fd_sc_hd__inv_2 _13473_ (.A(_09209_),
    .Y(_09210_));
 sky130_fd_sc_hd__nand3_1 _13474_ (.A(_09205_),
    .B(_09206_),
    .C(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_1 _13475_ (.A(_09211_),
    .B(_09206_),
    .Y(_09212_));
 sky130_fd_sc_hd__nand3_1 _13476_ (.A(_09199_),
    .B(_09147_),
    .C(_09143_),
    .Y(_09213_));
 sky130_fd_sc_hd__inv_2 _13477_ (.A(_09143_),
    .Y(_09214_));
 sky130_fd_sc_hd__nand2_1 _13478_ (.A(_09148_),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__nand2_1 _13479_ (.A(_09213_),
    .B(_09215_),
    .Y(_09216_));
 sky130_fd_sc_hd__nand2_1 _13480_ (.A(_09216_),
    .B(\base_h_sync[2] ),
    .Y(_09217_));
 sky130_fd_sc_hd__inv_2 _13481_ (.A(\base_h_sync[2] ),
    .Y(_09218_));
 sky130_fd_sc_hd__nand3_1 _13482_ (.A(_09213_),
    .B(_09218_),
    .C(_09215_),
    .Y(_09219_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(_09217_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__nand2_1 _13484_ (.A(_09212_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand3_1 _13485_ (.A(_09213_),
    .B(\base_h_sync[2] ),
    .C(_09215_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_1 _13486_ (.A(_09221_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__nand2_1 _13487_ (.A(_09215_),
    .B(_09142_),
    .Y(_09224_));
 sky130_fd_sc_hd__clkinvlp_2 _13488_ (.A(_09139_),
    .Y(_09225_));
 sky130_fd_sc_hd__nand2_1 _13489_ (.A(_09224_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__nand3_1 _13490_ (.A(_09215_),
    .B(_09139_),
    .C(_09142_),
    .Y(_09227_));
 sky130_fd_sc_hd__nand2_1 _13491_ (.A(_09226_),
    .B(_09227_),
    .Y(_09228_));
 sky130_fd_sc_hd__inv_2 _13492_ (.A(\base_h_sync[3] ),
    .Y(_09229_));
 sky130_fd_sc_hd__nand2_1 _13493_ (.A(_09228_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_1 _13494_ (.A(_09223_),
    .B(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__nand3_2 _13495_ (.A(_09226_),
    .B(\base_h_sync[3] ),
    .C(_09227_),
    .Y(_09232_));
 sky130_fd_sc_hd__nand2_1 _13496_ (.A(_09231_),
    .B(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__xor2_1 _13497_ (.A(\base_h_sync[4] ),
    .B(_09186_),
    .X(_09234_));
 sky130_fd_sc_hd__inv_2 _13498_ (.A(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand2_1 _13499_ (.A(_09182_),
    .B(\base_h_sync[5] ),
    .Y(_09236_));
 sky130_fd_sc_hd__nand3_1 _13500_ (.A(_09181_),
    .B(_09171_),
    .C(_09183_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_1 _13501_ (.A(_09236_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__nand2_1 _13502_ (.A(_09235_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__inv_2 _13503_ (.A(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__nand3_1 _13504_ (.A(_09179_),
    .B(_09233_),
    .C(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__inv_2 _13505_ (.A(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__nor2_1 _13506_ (.A(_09195_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__or2_1 _13507_ (.A(_09168_),
    .B(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__nand2_1 _13508_ (.A(_09243_),
    .B(_09168_),
    .Y(_09245_));
 sky130_fd_sc_hd__nand2_1 _13509_ (.A(_09244_),
    .B(_09245_),
    .Y(_09246_));
 sky130_fd_sc_hd__inv_2 _13510_ (.A(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__xor2_1 _13511_ (.A(\base_h_active[9] ),
    .B(_09167_),
    .X(_09248_));
 sky130_fd_sc_hd__inv_2 _13512_ (.A(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__xor2_2 _13513_ (.A(_09249_),
    .B(_09244_),
    .X(_09250_));
 sky130_fd_sc_hd__inv_2 _13514_ (.A(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__inv_2 _13515_ (.A(net3947),
    .Y(_09252_));
 sky130_fd_sc_hd__a22o_1 _13516_ (.A1(_08910_),
    .A2(_09247_),
    .B1(_09251_),
    .B2(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__nand3_1 _13517_ (.A(_09233_),
    .B(_09238_),
    .C(_09235_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand2_1 _13518_ (.A(_09254_),
    .B(_09191_),
    .Y(_09255_));
 sky130_fd_sc_hd__inv_2 _13519_ (.A(_09178_),
    .Y(_09256_));
 sky130_fd_sc_hd__nand2_1 _13520_ (.A(_09255_),
    .B(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__nand3_1 _13521_ (.A(_09257_),
    .B(_09170_),
    .C(_09177_),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_2 _13522_ (.A(_09258_),
    .B(_09243_),
    .Y(_09259_));
 sky130_fd_sc_hd__inv_2 _13523_ (.A(_09259_),
    .Y(_09260_));
 sky130_fd_sc_hd__nand2_1 _13524_ (.A(_09260_),
    .B(_08874_),
    .Y(_09261_));
 sky130_fd_sc_hd__nand2_2 _13525_ (.A(_09233_),
    .B(_09235_),
    .Y(_09262_));
 sky130_fd_sc_hd__nand2_1 _13526_ (.A(_09262_),
    .B(_09188_),
    .Y(_09263_));
 sky130_fd_sc_hd__nand2_1 _13527_ (.A(_09263_),
    .B(_09238_),
    .Y(_09264_));
 sky130_fd_sc_hd__inv_2 _13528_ (.A(_09238_),
    .Y(_09265_));
 sky130_fd_sc_hd__nand3_2 _13529_ (.A(_09262_),
    .B(_09265_),
    .C(_09188_),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_1 _13530_ (.A(_09264_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__nand3_1 _13531_ (.A(_09231_),
    .B(_09234_),
    .C(_09232_),
    .Y(_09268_));
 sky130_fd_sc_hd__nand2_1 _13532_ (.A(_09262_),
    .B(_09268_),
    .Y(_09269_));
 sky130_fd_sc_hd__nand2_1 _13533_ (.A(_09216_),
    .B(_09218_),
    .Y(_09270_));
 sky130_fd_sc_hd__nand2_1 _13534_ (.A(_09270_),
    .B(_09222_),
    .Y(_09271_));
 sky130_fd_sc_hd__a21boi_1 _13535_ (.A1(_09205_),
    .A2(_09210_),
    .B1_N(_09206_),
    .Y(_09272_));
 sky130_fd_sc_hd__nand2_1 _13536_ (.A(_09271_),
    .B(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_1 _13537_ (.A(_09221_),
    .B(_09273_),
    .Y(_09274_));
 sky130_fd_sc_hd__nand3_1 _13538_ (.A(_09223_),
    .B(_09232_),
    .C(_09230_),
    .Y(_09275_));
 sky130_fd_sc_hd__nand2_1 _13539_ (.A(_09230_),
    .B(_09232_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand3_1 _13540_ (.A(_09276_),
    .B(_09222_),
    .C(_09221_),
    .Y(_09277_));
 sky130_fd_sc_hd__nand2_1 _13541_ (.A(_09275_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_09203_),
    .B(\base_h_sync[1] ),
    .Y(_09279_));
 sky130_fd_sc_hd__nand3_1 _13543_ (.A(_09199_),
    .B(_09202_),
    .C(_09204_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand3_1 _13544_ (.A(_09279_),
    .B(_09280_),
    .C(_09209_),
    .Y(_09281_));
 sky130_fd_sc_hd__nand2_1 _13545_ (.A(_09211_),
    .B(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__nand2_1 _13546_ (.A(_09282_),
    .B(\base_h_counter[1] ),
    .Y(_09283_));
 sky130_fd_sc_hd__or2_1 _13547_ (.A(\base_h_sync[0] ),
    .B(_09208_),
    .X(_09284_));
 sky130_fd_sc_hd__nand2_1 _13548_ (.A(_09284_),
    .B(_09209_),
    .Y(_09285_));
 sky130_fd_sc_hd__inv_2 _13549_ (.A(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__nor2_1 _13550_ (.A(\base_h_counter[1] ),
    .B(_09282_),
    .Y(_09287_));
 sky130_fd_sc_hd__a31o_1 _13551_ (.A1(_09283_),
    .A2(_08890_),
    .A3(_09286_),
    .B1(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__nand2_1 _13552_ (.A(_09274_),
    .B(\base_h_counter[2] ),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_1 _13553_ (.A(_09288_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__o221ai_1 _13554_ (.A1(\base_h_counter[2] ),
    .A2(_09274_),
    .B1(\base_h_counter[3] ),
    .B2(_09278_),
    .C1(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__nand2_1 _13555_ (.A(_09269_),
    .B(\base_h_counter[4] ),
    .Y(_09292_));
 sky130_fd_sc_hd__nand2_1 _13556_ (.A(_09278_),
    .B(\base_h_counter[3] ),
    .Y(_09293_));
 sky130_fd_sc_hd__nand3_1 _13557_ (.A(_09291_),
    .B(_09292_),
    .C(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__o221ai_1 _13558_ (.A1(\base_h_counter[5] ),
    .A2(_09267_),
    .B1(\base_h_counter[4] ),
    .B2(_09269_),
    .C1(_09294_),
    .Y(_09295_));
 sky130_fd_sc_hd__nand3_1 _13559_ (.A(_09254_),
    .B(_09178_),
    .C(_09191_),
    .Y(_09296_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(_09257_),
    .B(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_1 _13561_ (.A(_09297_),
    .B(\base_h_counter[6] ),
    .Y(_09298_));
 sky130_fd_sc_hd__nand2_1 _13562_ (.A(_09267_),
    .B(\base_h_counter[5] ),
    .Y(_09299_));
 sky130_fd_sc_hd__nand3_1 _13563_ (.A(_09295_),
    .B(_09298_),
    .C(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__or2_1 _13564_ (.A(\base_h_counter[6] ),
    .B(_09297_),
    .X(_09301_));
 sky130_fd_sc_hd__a22o_1 _13565_ (.A1(\base_h_counter[7] ),
    .A2(_09259_),
    .B1(_09300_),
    .B2(_09301_),
    .X(_09302_));
 sky130_fd_sc_hd__o2bb2a_1 _13566_ (.A1_N(_09261_),
    .A2_N(_09302_),
    .B1(_08910_),
    .B2(_09247_),
    .X(_09303_));
 sky130_fd_sc_hd__nand2_1 _13567_ (.A(_09250_),
    .B(\base_h_counter[9] ),
    .Y(_09304_));
 sky130_fd_sc_hd__or2_1 _13568_ (.A(\base_h_counter[8] ),
    .B(_09168_),
    .X(_09305_));
 sky130_fd_sc_hd__inv_2 _13569_ (.A(_09170_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_1 _13570_ (.A(_09228_),
    .B(\base_h_counter[3] ),
    .Y(_09307_));
 sky130_fd_sc_hd__nand2_1 _13571_ (.A(_09186_),
    .B(\base_h_counter[4] ),
    .Y(_09308_));
 sky130_fd_sc_hd__nand2_1 _13572_ (.A(_09187_),
    .B(_08879_),
    .Y(_09309_));
 sky130_fd_sc_hd__o21ai_1 _13573_ (.A1(\base_h_counter[5] ),
    .A2(_09182_),
    .B1(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__a21o_1 _13574_ (.A1(_09307_),
    .A2(_09308_),
    .B1(_09310_),
    .X(_09311_));
 sky130_fd_sc_hd__and2_1 _13575_ (.A(_09216_),
    .B(\base_h_counter[2] ),
    .X(_09312_));
 sky130_fd_sc_hd__nand2_1 _13576_ (.A(_09203_),
    .B(\base_h_counter[1] ),
    .Y(_09313_));
 sky130_fd_sc_hd__and3_1 _13577_ (.A(_09313_),
    .B(_08890_),
    .C(_09208_),
    .X(_09314_));
 sky130_fd_sc_hd__o21ba_1 _13578_ (.A1(\base_h_counter[1] ),
    .A2(_09203_),
    .B1_N(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__or2_1 _13579_ (.A(\base_h_counter[3] ),
    .B(_09228_),
    .X(_09316_));
 sky130_fd_sc_hd__or2_1 _13580_ (.A(\base_h_counter[2] ),
    .B(_09216_),
    .X(_09317_));
 sky130_fd_sc_hd__o211ai_1 _13581_ (.A1(_09312_),
    .A2(_09315_),
    .B1(_09316_),
    .C1(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__nand2_1 _13582_ (.A(_09182_),
    .B(\base_h_counter[5] ),
    .Y(_09319_));
 sky130_fd_sc_hd__nand2_1 _13583_ (.A(_09174_),
    .B(\base_h_counter[6] ),
    .Y(_09320_));
 sky130_fd_sc_hd__o211a_1 _13584_ (.A1(_09310_),
    .A2(_09318_),
    .B1(_09319_),
    .C1(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__a2bb2o_1 _13585_ (.A1_N(\base_h_counter[6] ),
    .A2_N(_09174_),
    .B1(_09311_),
    .B2(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__o21ai_1 _13586_ (.A1(_08874_),
    .A2(_09306_),
    .B1(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__nand2_1 _13587_ (.A(_09306_),
    .B(_08874_),
    .Y(_09324_));
 sky130_fd_sc_hd__a22o_1 _13588_ (.A1(\base_h_counter[8] ),
    .A2(_09168_),
    .B1(_09323_),
    .B2(_09324_),
    .X(_09325_));
 sky130_fd_sc_hd__o211ai_1 _13589_ (.A1(\base_h_counter[9] ),
    .A2(_09248_),
    .B1(_09305_),
    .C1(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__o21ai_1 _13590_ (.A1(_09252_),
    .A2(_09249_),
    .B1(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__o211a_4 _13591_ (.A1(_09253_),
    .A2(_09303_),
    .B1(_09304_),
    .C1(_09327_),
    .X(net92));
 sky130_fd_sc_hd__or2_1 _13592_ (.A(\base_v_active[0] ),
    .B(\base_v_fporch[0] ),
    .X(_09328_));
 sky130_fd_sc_hd__nand2_1 _13593_ (.A(\base_v_active[0] ),
    .B(\base_v_fporch[0] ),
    .Y(_09329_));
 sky130_fd_sc_hd__nand2_1 _13594_ (.A(_09328_),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__inv_2 _13595_ (.A(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__inv_2 _13596_ (.A(\base_v_fporch[1] ),
    .Y(_09332_));
 sky130_fd_sc_hd__nand2_1 _13597_ (.A(_08953_),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_1 _13598_ (.A(\base_v_active[1] ),
    .B(\base_v_fporch[1] ),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _13599_ (.A(_09333_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__or2_1 _13600_ (.A(_09329_),
    .B(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__nand2_1 _13601_ (.A(_09335_),
    .B(_09329_),
    .Y(_09337_));
 sky130_fd_sc_hd__nand2_1 _13602_ (.A(_09336_),
    .B(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__inv_2 _13603_ (.A(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__inv_2 _13604_ (.A(net3800),
    .Y(_09340_));
 sky130_fd_sc_hd__nand2_1 _13605_ (.A(_09339_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__o21ai_1 _13606_ (.A1(_08938_),
    .A2(_09331_),
    .B1(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__a21o_1 _13607_ (.A1(\base_v_counter[1] ),
    .A2(_09338_),
    .B1(_09342_),
    .X(_09343_));
 sky130_fd_sc_hd__nand2_1 _13608_ (.A(_09336_),
    .B(_09334_),
    .Y(_09344_));
 sky130_fd_sc_hd__or2_1 _13609_ (.A(\base_v_active[2] ),
    .B(\base_v_fporch[2] ),
    .X(_09345_));
 sky130_fd_sc_hd__nand2_1 _13610_ (.A(\base_v_active[2] ),
    .B(\base_v_fporch[2] ),
    .Y(_09346_));
 sky130_fd_sc_hd__nand2_1 _13611_ (.A(_09345_),
    .B(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__inv_2 _13612_ (.A(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__nand2_1 _13613_ (.A(_09344_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__and2_1 _13614_ (.A(_09349_),
    .B(_09346_),
    .X(_09350_));
 sky130_fd_sc_hd__or2_1 _13615_ (.A(_08946_),
    .B(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__nand2_1 _13616_ (.A(_09350_),
    .B(_08946_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_1 _13617_ (.A(_09351_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__nor2_1 _13618_ (.A(\base_v_counter[3] ),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__inv_2 _13619_ (.A(_09353_),
    .Y(_09355_));
 sky130_fd_sc_hd__nor2_1 _13620_ (.A(_08944_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__nor2_1 _13621_ (.A(_09354_),
    .B(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__or2_1 _13622_ (.A(_09348_),
    .B(_09344_),
    .X(_09358_));
 sky130_fd_sc_hd__nand2_1 _13623_ (.A(_09358_),
    .B(_09349_),
    .Y(_09359_));
 sky130_fd_sc_hd__inv_2 _13624_ (.A(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__nand2_1 _13625_ (.A(_09360_),
    .B(_08949_),
    .Y(_09361_));
 sky130_fd_sc_hd__nand2_1 _13626_ (.A(_09359_),
    .B(\base_v_counter[2] ),
    .Y(_09362_));
 sky130_fd_sc_hd__nand3_1 _13627_ (.A(_09357_),
    .B(_09361_),
    .C(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__a211o_1 _13628_ (.A1(_08938_),
    .A2(_09331_),
    .B1(_09343_),
    .C1(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__nand3b_2 _13629_ (.A_N(_09350_),
    .B(\base_v_active[4] ),
    .C(\base_v_active[3] ),
    .Y(_09365_));
 sky130_fd_sc_hd__nor2_1 _13630_ (.A(_08927_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__inv_2 _13631_ (.A(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand2_1 _13632_ (.A(_09365_),
    .B(_08927_),
    .Y(_09368_));
 sky130_fd_sc_hd__nand2_1 _13633_ (.A(_09367_),
    .B(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__inv_2 _13634_ (.A(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__nand2_1 _13635_ (.A(_09370_),
    .B(_08929_),
    .Y(_09371_));
 sky130_fd_sc_hd__nand2_1 _13636_ (.A(_09369_),
    .B(\base_v_counter[5] ),
    .Y(_09372_));
 sky130_fd_sc_hd__nand2_1 _13637_ (.A(_09371_),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_1 _13638_ (.A(_09351_),
    .B(_08932_),
    .Y(_09374_));
 sky130_fd_sc_hd__nand2_1 _13639_ (.A(_09374_),
    .B(_09365_),
    .Y(_09375_));
 sky130_fd_sc_hd__or2_1 _13640_ (.A(\base_v_counter[4] ),
    .B(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__nand2_1 _13641_ (.A(_09375_),
    .B(\base_v_counter[4] ),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_1 _13642_ (.A(_09376_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__nand2_1 _13643_ (.A(_09367_),
    .B(_08915_),
    .Y(_09379_));
 sky130_fd_sc_hd__nand2_1 _13644_ (.A(_09366_),
    .B(\base_v_active[6] ),
    .Y(_09380_));
 sky130_fd_sc_hd__nand2_1 _13645_ (.A(_09379_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__inv_2 _13646_ (.A(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__nor2_1 _13647_ (.A(_08917_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand2_1 _13648_ (.A(_09380_),
    .B(_08922_),
    .Y(_09384_));
 sky130_fd_sc_hd__nand3_1 _13649_ (.A(_09366_),
    .B(\base_v_active[7] ),
    .C(\base_v_active[6] ),
    .Y(_09385_));
 sky130_fd_sc_hd__nand2_1 _13650_ (.A(_09384_),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__xor2_1 _13651_ (.A(_08919_),
    .B(_09386_),
    .X(_09387_));
 sky130_fd_sc_hd__inv_2 _13652_ (.A(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(_09382_),
    .B(_08917_),
    .Y(_09389_));
 sky130_fd_sc_hd__or3b_1 _13654_ (.A(_09383_),
    .B(_09388_),
    .C_N(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__nor3_1 _13655_ (.A(_09373_),
    .B(_09378_),
    .C(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__or2_1 _13656_ (.A(_08939_),
    .B(_09385_),
    .X(_09392_));
 sky130_fd_sc_hd__buf_6 _13657_ (.A(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__xor2_1 _13658_ (.A(\base_v_counter[9] ),
    .B(_09393_),
    .X(_09394_));
 sky130_fd_sc_hd__nand2_1 _13659_ (.A(_09385_),
    .B(_08939_),
    .Y(_09395_));
 sky130_fd_sc_hd__nand2_1 _13660_ (.A(_09393_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__inv_2 _13661_ (.A(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__nand2_1 _13662_ (.A(_09397_),
    .B(_08941_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand2_1 _13663_ (.A(_09396_),
    .B(\base_v_counter[8] ),
    .Y(_09399_));
 sky130_fd_sc_hd__and3_1 _13664_ (.A(_09394_),
    .B(_09398_),
    .C(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__and3b_1 _13665_ (.A_N(_09364_),
    .B(_09391_),
    .C(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__o21a_1 _13666_ (.A1(_09376_),
    .A2(_09373_),
    .B1(_09371_),
    .X(_09402_));
 sky130_fd_sc_hd__inv_2 _13667_ (.A(_09386_),
    .Y(_09403_));
 sky130_fd_sc_hd__nand2_1 _13668_ (.A(_09403_),
    .B(_08920_),
    .Y(_09404_));
 sky130_fd_sc_hd__o221a_1 _13669_ (.A1(_09389_),
    .A2(_09388_),
    .B1(_09402_),
    .B2(_09390_),
    .C1(_09404_),
    .X(_09405_));
 sky130_fd_sc_hd__a21oi_1 _13670_ (.A1(_09341_),
    .A2(_09343_),
    .B1(_09363_),
    .Y(_09406_));
 sky130_fd_sc_hd__a311o_1 _13671_ (.A1(_08949_),
    .A2(_09360_),
    .A3(_09357_),
    .B1(_09354_),
    .C1(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__nand2_1 _13672_ (.A(_09391_),
    .B(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_1 _13673_ (.A(_09405_),
    .B(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__nor2_1 _13674_ (.A(\base_v_counter[9] ),
    .B(_09393_),
    .Y(_09410_));
 sky130_fd_sc_hd__a31o_1 _13675_ (.A1(_09394_),
    .A2(_08941_),
    .A3(_09397_),
    .B1(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__a21oi_1 _13676_ (.A1(_09409_),
    .A2(_09400_),
    .B1(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__nand2_1 _13677_ (.A(_09339_),
    .B(\base_v_sync[1] ),
    .Y(_09413_));
 sky130_fd_sc_hd__nand2_1 _13678_ (.A(_09331_),
    .B(\base_v_sync[0] ),
    .Y(_09414_));
 sky130_fd_sc_hd__inv_2 _13679_ (.A(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__inv_2 _13680_ (.A(\base_v_sync[1] ),
    .Y(_09416_));
 sky130_fd_sc_hd__nand2_1 _13681_ (.A(_09338_),
    .B(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__nand3_1 _13682_ (.A(_09413_),
    .B(_09415_),
    .C(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__nand2_1 _13683_ (.A(_09418_),
    .B(_09413_),
    .Y(_09419_));
 sky130_fd_sc_hd__inv_2 _13684_ (.A(\base_v_sync[2] ),
    .Y(_09420_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(_09359_),
    .B(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand3_2 _13686_ (.A(_09358_),
    .B(\base_v_sync[2] ),
    .C(_09349_),
    .Y(_09422_));
 sky130_fd_sc_hd__nand3_2 _13687_ (.A(_09419_),
    .B(_09421_),
    .C(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__nand2_1 _13688_ (.A(_09423_),
    .B(_09422_),
    .Y(_09424_));
 sky130_fd_sc_hd__nand2_1 _13689_ (.A(_09424_),
    .B(_09355_),
    .Y(_09425_));
 sky130_fd_sc_hd__or2_1 _13690_ (.A(_09375_),
    .B(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__nand2_1 _13691_ (.A(_09425_),
    .B(_09375_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_1 _13692_ (.A(_09426_),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__inv_2 _13693_ (.A(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__nor2_1 _13694_ (.A(_08934_),
    .B(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__nor2_1 _13695_ (.A(\base_v_counter[4] ),
    .B(_09428_),
    .Y(_09431_));
 sky130_fd_sc_hd__nand2_1 _13696_ (.A(_09426_),
    .B(_09369_),
    .Y(_09432_));
 sky130_fd_sc_hd__nand3_1 _13697_ (.A(_09374_),
    .B(\base_v_active[5] ),
    .C(_09365_),
    .Y(_09433_));
 sky130_fd_sc_hd__or2_1 _13698_ (.A(_09433_),
    .B(_09425_),
    .X(_09434_));
 sky130_fd_sc_hd__nand2_1 _13699_ (.A(_09432_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__or2_1 _13700_ (.A(\base_v_counter[5] ),
    .B(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__nand2_1 _13701_ (.A(_09435_),
    .B(\base_v_counter[5] ),
    .Y(_09437_));
 sky130_fd_sc_hd__nand2_1 _13702_ (.A(_09436_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__or3_1 _13703_ (.A(_09430_),
    .B(_09431_),
    .C(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__nor2_1 _13704_ (.A(_09381_),
    .B(_09434_),
    .Y(_09440_));
 sky130_fd_sc_hd__inv_2 _13705_ (.A(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__nand2_1 _13706_ (.A(_09441_),
    .B(_09386_),
    .Y(_09442_));
 sky130_fd_sc_hd__nand2_1 _13707_ (.A(_09440_),
    .B(_09403_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand2_1 _13708_ (.A(_09442_),
    .B(_09443_),
    .Y(_09444_));
 sky130_fd_sc_hd__xor2_1 _13709_ (.A(_08919_),
    .B(_09444_),
    .X(_09445_));
 sky130_fd_sc_hd__nand2_1 _13710_ (.A(_09434_),
    .B(_09381_),
    .Y(_09446_));
 sky130_fd_sc_hd__nand2_1 _13711_ (.A(_09441_),
    .B(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__nor2_1 _13712_ (.A(\base_v_counter[6] ),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__inv_2 _13713_ (.A(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nand2_1 _13714_ (.A(_09447_),
    .B(\base_v_counter[6] ),
    .Y(_09450_));
 sky130_fd_sc_hd__and3_1 _13715_ (.A(_09445_),
    .B(_09449_),
    .C(_09450_),
    .X(_09451_));
 sky130_fd_sc_hd__and2b_1 _13716_ (.A_N(_09439_),
    .B(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__or2_1 _13717_ (.A(_09396_),
    .B(_09443_),
    .X(_09453_));
 sky130_fd_sc_hd__nand2_1 _13718_ (.A(_09453_),
    .B(_09393_),
    .Y(_09454_));
 sky130_fd_sc_hd__xor2_1 _13719_ (.A(_08960_),
    .B(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__nand2_1 _13720_ (.A(_09443_),
    .B(_09396_),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_1 _13721_ (.A(_09453_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__inv_2 _13722_ (.A(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__nand2_1 _13723_ (.A(_09458_),
    .B(_08941_),
    .Y(_09459_));
 sky130_fd_sc_hd__nand2_1 _13724_ (.A(_09457_),
    .B(\base_v_counter[8] ),
    .Y(_09460_));
 sky130_fd_sc_hd__and3_1 _13725_ (.A(_09455_),
    .B(_09459_),
    .C(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__or2_1 _13726_ (.A(\base_v_sync[0] ),
    .B(_09331_),
    .X(_09462_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(_09462_),
    .B(_09414_),
    .Y(_09463_));
 sky130_fd_sc_hd__inv_2 _13728_ (.A(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand2_1 _13729_ (.A(_09413_),
    .B(_09417_),
    .Y(_09465_));
 sky130_fd_sc_hd__nand2_1 _13730_ (.A(_09465_),
    .B(_09414_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand2_1 _13731_ (.A(_09466_),
    .B(_09418_),
    .Y(_09467_));
 sky130_fd_sc_hd__nand2_1 _13732_ (.A(_09467_),
    .B(\base_v_counter[1] ),
    .Y(_09468_));
 sky130_fd_sc_hd__or2_1 _13733_ (.A(\base_v_counter[1] ),
    .B(_09467_),
    .X(_09469_));
 sky130_fd_sc_hd__o211ai_1 _13734_ (.A1(_08938_),
    .A2(_09464_),
    .B1(_09468_),
    .C1(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__nand3_1 _13735_ (.A(_09423_),
    .B(_09353_),
    .C(_09422_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand2_1 _13736_ (.A(_09425_),
    .B(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__or2_1 _13737_ (.A(\base_v_counter[3] ),
    .B(_09472_),
    .X(_09473_));
 sky130_fd_sc_hd__a21o_1 _13738_ (.A1(_09421_),
    .A2(_09422_),
    .B1(_09419_),
    .X(_09474_));
 sky130_fd_sc_hd__nand2_1 _13739_ (.A(_09474_),
    .B(_09423_),
    .Y(_09475_));
 sky130_fd_sc_hd__or2_1 _13740_ (.A(\base_v_counter[2] ),
    .B(_09475_),
    .X(_09476_));
 sky130_fd_sc_hd__nand2_1 _13741_ (.A(_09475_),
    .B(\base_v_counter[2] ),
    .Y(_09477_));
 sky130_fd_sc_hd__nand2_1 _13742_ (.A(_09472_),
    .B(\base_v_counter[3] ),
    .Y(_09478_));
 sky130_fd_sc_hd__and4_1 _13743_ (.A(_09473_),
    .B(_09476_),
    .C(_09477_),
    .D(_09478_),
    .X(_09479_));
 sky130_fd_sc_hd__inv_2 _13744_ (.A(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__a211oi_1 _13745_ (.A1(_08938_),
    .A2(_09464_),
    .B1(_09470_),
    .C1(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__nand3_1 _13746_ (.A(_09452_),
    .B(_09461_),
    .C(_09481_),
    .Y(_09482_));
 sky130_fd_sc_hd__nand2_1 _13747_ (.A(_09473_),
    .B(_09478_),
    .Y(_09483_));
 sky130_fd_sc_hd__and2_1 _13748_ (.A(_09470_),
    .B(_09469_),
    .X(_09484_));
 sky130_fd_sc_hd__o221ai_2 _13749_ (.A1(_09476_),
    .A2(_09483_),
    .B1(_09484_),
    .B2(_09480_),
    .C1(_09473_),
    .Y(_09485_));
 sky130_fd_sc_hd__nand2_1 _13750_ (.A(_09445_),
    .B(_09448_),
    .Y(_09486_));
 sky130_fd_sc_hd__a21bo_1 _13751_ (.A1(_09431_),
    .A2(_09437_),
    .B1_N(_09436_),
    .X(_09487_));
 sky130_fd_sc_hd__nand2_1 _13752_ (.A(_09451_),
    .B(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__o211ai_1 _13753_ (.A1(_08919_),
    .A2(_09444_),
    .B1(_09486_),
    .C1(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__a21o_1 _13754_ (.A1(_09485_),
    .A2(_09452_),
    .B1(_09489_),
    .X(_09490_));
 sky130_fd_sc_hd__inv_2 _13755_ (.A(_09454_),
    .Y(_09491_));
 sky130_fd_sc_hd__nor2_1 _13756_ (.A(\base_v_counter[9] ),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__a31o_1 _13757_ (.A1(_09455_),
    .A2(_08941_),
    .A3(_09458_),
    .B1(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__a21o_1 _13758_ (.A1(_09490_),
    .A2(_09461_),
    .B1(_09493_),
    .X(_09494_));
 sky130_fd_sc_hd__o211ai_4 _13759_ (.A1(_09401_),
    .A2(_09412_),
    .B1(_09482_),
    .C1(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__inv_2 _13760_ (.A(net135),
    .Y(net134));
 sky130_fd_sc_hd__nand2_2 _13761_ (.A(_08848_),
    .B(_09125_),
    .Y(_09496_));
 sky130_fd_sc_hd__clkbuf_8 _13762_ (.A(_09496_),
    .X(_09497_));
 sky130_fd_sc_hd__inv_2 _13763_ (.A(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_1 _13764_ (.A(_09498_),
    .B(_08840_),
    .Y(_09499_));
 sky130_fd_sc_hd__inv_2 _13765_ (.A(_09499_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _13766_ (.A(net2387),
    .B(net3958),
    .Y(_09500_));
 sky130_fd_sc_hd__nand2_1 _13767_ (.A(net2387),
    .B(net3958),
    .Y(_09501_));
 sky130_fd_sc_hd__inv_2 _13768_ (.A(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__or3_1 _13769_ (.A(_09500_),
    .B(_09502_),
    .C(_09497_),
    .X(_09503_));
 sky130_fd_sc_hd__inv_2 _13770_ (.A(_09503_),
    .Y(_00001_));
 sky130_fd_sc_hd__inv_2 _13771_ (.A(net3991),
    .Y(_09504_));
 sky130_fd_sc_hd__nor2_1 _13772_ (.A(_09504_),
    .B(_09501_),
    .Y(_09505_));
 sky130_fd_sc_hd__nor2_1 _13773_ (.A(net3991),
    .B(_09502_),
    .Y(_09506_));
 sky130_fd_sc_hd__or3_1 _13774_ (.A(_09505_),
    .B(_09506_),
    .C(_09497_),
    .X(_09507_));
 sky130_fd_sc_hd__inv_2 _13775_ (.A(_09507_),
    .Y(_00002_));
 sky130_fd_sc_hd__and2_1 _13776_ (.A(_09505_),
    .B(net4000),
    .X(_09508_));
 sky130_fd_sc_hd__or2_1 _13777_ (.A(net4000),
    .B(_09505_),
    .X(_09509_));
 sky130_fd_sc_hd__or3b_1 _13778_ (.A(_09508_),
    .B(_09497_),
    .C_N(_09509_),
    .X(_09510_));
 sky130_fd_sc_hd__inv_2 _13779_ (.A(_09510_),
    .Y(_00003_));
 sky130_fd_sc_hd__nor2_1 _13780_ (.A(net3984),
    .B(_09508_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_1 _13781_ (.A(_09508_),
    .B(net3984),
    .Y(_09512_));
 sky130_fd_sc_hd__or3b_1 _13782_ (.A(_09130_),
    .B(net3985),
    .C_N(_09512_),
    .X(_09513_));
 sky130_fd_sc_hd__inv_2 _13783_ (.A(net3986),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _13784_ (.A(net3888),
    .Y(_09514_));
 sky130_fd_sc_hd__or2_1 _13785_ (.A(_09514_),
    .B(_09512_),
    .X(_09515_));
 sky130_fd_sc_hd__buf_6 _13786_ (.A(_09126_),
    .X(_09516_));
 sky130_fd_sc_hd__nand2_1 _13787_ (.A(_09512_),
    .B(_09514_),
    .Y(_09517_));
 sky130_fd_sc_hd__nand3_1 _13788_ (.A(_09515_),
    .B(_09516_),
    .C(net3889),
    .Y(_09518_));
 sky130_fd_sc_hd__inv_2 _13789_ (.A(net3890),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_2 _13790_ (.A(net3872),
    .Y(_09519_));
 sky130_fd_sc_hd__or2_1 _13791_ (.A(_09519_),
    .B(_09515_),
    .X(_09520_));
 sky130_fd_sc_hd__nand2_1 _13792_ (.A(_09515_),
    .B(_09519_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand3_1 _13793_ (.A(_09520_),
    .B(_09516_),
    .C(net3873),
    .Y(_09522_));
 sky130_fd_sc_hd__inv_2 _13794_ (.A(net3874),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_2 _13795_ (.A(net3997),
    .Y(_09523_));
 sky130_fd_sc_hd__nor2_1 _13796_ (.A(_09523_),
    .B(_09520_),
    .Y(_09524_));
 sky130_fd_sc_hd__nand2_1 _13797_ (.A(_09520_),
    .B(_09523_),
    .Y(_09525_));
 sky130_fd_sc_hd__or3b_1 _13798_ (.A(_09130_),
    .B(_09524_),
    .C_N(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__inv_2 _13799_ (.A(_09526_),
    .Y(_00007_));
 sky130_fd_sc_hd__or2_1 _13800_ (.A(net3979),
    .B(_09524_),
    .X(_09527_));
 sky130_fd_sc_hd__nand2_1 _13801_ (.A(_09524_),
    .B(net3979),
    .Y(_09528_));
 sky130_fd_sc_hd__and3_1 _13802_ (.A(net3980),
    .B(_09516_),
    .C(_09528_),
    .X(_09529_));
 sky130_fd_sc_hd__clkbuf_1 _13803_ (.A(net3981),
    .X(_00008_));
 sky130_fd_sc_hd__buf_8 _13804_ (.A(_08995_),
    .X(_09530_));
 sky130_fd_sc_hd__clkbuf_16 _13805_ (.A(_09530_),
    .X(_09531_));
 sky130_fd_sc_hd__buf_6 _13806_ (.A(_09531_),
    .X(_09532_));
 sky130_fd_sc_hd__clkbuf_8 _13807_ (.A(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(\res_h_counter[6] ),
    .B(\res_h_counter[7] ),
    .Y(_09534_));
 sky130_fd_sc_hd__inv_6 _13809_ (.A(_09534_),
    .Y(_09535_));
 sky130_fd_sc_hd__nor2_8 _13810_ (.A(\res_h_counter[4] ),
    .B(\res_h_counter[5] ),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_8 _13811_ (.A(_09535_),
    .B(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__inv_2 _13812_ (.A(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__clkbuf_4 _13813_ (.A(_09538_),
    .X(_09539_));
 sky130_fd_sc_hd__clkbuf_4 _13814_ (.A(_09539_),
    .X(_09540_));
 sky130_fd_sc_hd__buf_12 _13815_ (.A(_08993_),
    .X(_09541_));
 sky130_fd_sc_hd__nor2_4 _13816_ (.A(\res_h_counter[5] ),
    .B(_09047_),
    .Y(_09542_));
 sky130_fd_sc_hd__nand2_8 _13817_ (.A(_09542_),
    .B(_09535_),
    .Y(_09543_));
 sky130_fd_sc_hd__nor2_4 _13818_ (.A(_09541_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__buf_8 _13819_ (.A(_09541_),
    .X(_09545_));
 sky130_fd_sc_hd__buf_6 _13820_ (.A(_09545_),
    .X(_09546_));
 sky130_fd_sc_hd__buf_6 _13821_ (.A(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__buf_8 _13822_ (.A(_09547_),
    .X(_09548_));
 sky130_fd_sc_hd__nor2_8 _13823_ (.A(\res_h_counter[4] ),
    .B(_09043_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2_8 _13824_ (.A(_09549_),
    .B(_09535_),
    .Y(_09550_));
 sky130_fd_sc_hd__buf_4 _13825_ (.A(_09541_),
    .X(_09551_));
 sky130_fd_sc_hd__nand2_1 _13826_ (.A(\res_h_counter[4] ),
    .B(\res_h_counter[5] ),
    .Y(_09552_));
 sky130_fd_sc_hd__clkinv_4 _13827_ (.A(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__nand2_8 _13828_ (.A(_09553_),
    .B(_09535_),
    .Y(_09554_));
 sky130_fd_sc_hd__buf_6 _13829_ (.A(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__and2_4 _13830_ (.A(_09017_),
    .B(net3867),
    .X(_09556_));
 sky130_fd_sc_hd__nor2_2 _13831_ (.A(\res_h_counter[2] ),
    .B(\res_h_counter[3] ),
    .Y(_09557_));
 sky130_fd_sc_hd__and2_4 _13832_ (.A(_09556_),
    .B(_09557_),
    .X(_09558_));
 sky130_fd_sc_hd__inv_2 _13833_ (.A(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__or3_1 _13834_ (.A(_09551_),
    .B(_09555_),
    .C(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__nand2_2 _13835_ (.A(\res_h_counter[0] ),
    .B(\res_h_counter[1] ),
    .Y(_09561_));
 sky130_fd_sc_hd__inv_2 _13836_ (.A(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__and2_4 _13837_ (.A(_09562_),
    .B(_09557_),
    .X(_09563_));
 sky130_fd_sc_hd__inv_2 _13838_ (.A(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__or3_1 _13839_ (.A(_09551_),
    .B(_09554_),
    .C(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__nor2_4 _13840_ (.A(net3867),
    .B(_09017_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand2_2 _13841_ (.A(_09566_),
    .B(_09557_),
    .Y(_09567_));
 sky130_fd_sc_hd__clkinv_4 _13842_ (.A(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__nand2_8 _13843_ (.A(_09568_),
    .B(_08995_),
    .Y(_09569_));
 sky130_fd_sc_hd__or2_4 _13844_ (.A(_09554_),
    .B(_09569_),
    .X(_09570_));
 sky130_fd_sc_hd__nor2_4 _13845_ (.A(\res_h_counter[0] ),
    .B(\res_h_counter[1] ),
    .Y(_09571_));
 sky130_fd_sc_hd__nand2_2 _13846_ (.A(_09571_),
    .B(_09557_),
    .Y(_09572_));
 sky130_fd_sc_hd__or3_1 _13847_ (.A(_09551_),
    .B(_09572_),
    .C(_09554_),
    .X(_09573_));
 sky130_fd_sc_hd__and4_1 _13848_ (.A(_09560_),
    .B(_09565_),
    .C(_09570_),
    .D(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__nor2_4 _13849_ (.A(\res_h_counter[2] ),
    .B(_09021_),
    .Y(_09575_));
 sky130_fd_sc_hd__nand2_2 _13850_ (.A(_09575_),
    .B(_09571_),
    .Y(_09576_));
 sky130_fd_sc_hd__inv_6 _13851_ (.A(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__nand2_8 _13852_ (.A(_09577_),
    .B(_08995_),
    .Y(_09578_));
 sky130_fd_sc_hd__nand2_4 _13853_ (.A(_09575_),
    .B(_09566_),
    .Y(_09579_));
 sky130_fd_sc_hd__or3_1 _13854_ (.A(_09551_),
    .B(_09555_),
    .C(_09579_),
    .X(_09580_));
 sky130_fd_sc_hd__nand2_4 _13855_ (.A(_09556_),
    .B(_09575_),
    .Y(_09581_));
 sky130_fd_sc_hd__or3_1 _13856_ (.A(_09551_),
    .B(_09555_),
    .C(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__clkbuf_8 _13857_ (.A(_09541_),
    .X(_09583_));
 sky130_fd_sc_hd__nand2_4 _13858_ (.A(_09575_),
    .B(_09562_),
    .Y(_09584_));
 sky130_fd_sc_hd__or3_1 _13859_ (.A(_09583_),
    .B(_09555_),
    .C(_09584_),
    .X(_09585_));
 sky130_fd_sc_hd__o2111a_1 _13860_ (.A1(_09555_),
    .A2(_09578_),
    .B1(_09580_),
    .C1(_09582_),
    .D1(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__nor2_4 _13861_ (.A(\res_h_counter[3] ),
    .B(_09029_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand2_4 _13862_ (.A(_09587_),
    .B(_09571_),
    .Y(_09588_));
 sky130_fd_sc_hd__or3_1 _13863_ (.A(_09551_),
    .B(_09554_),
    .C(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_4 _13864_ (.A(_09556_),
    .B(_09587_),
    .Y(_09590_));
 sky130_fd_sc_hd__or3_1 _13865_ (.A(_09545_),
    .B(_09554_),
    .C(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__nand2_4 _13866_ (.A(_09587_),
    .B(_09562_),
    .Y(_09592_));
 sky130_fd_sc_hd__or3_1 _13867_ (.A(_09545_),
    .B(_09554_),
    .C(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__nand2_4 _13868_ (.A(_09587_),
    .B(_09566_),
    .Y(_09594_));
 sky130_fd_sc_hd__nor2_8 _13869_ (.A(_08993_),
    .B(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__inv_12 _13870_ (.A(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__or2_4 _13871_ (.A(_09554_),
    .B(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__and4_1 _13872_ (.A(_09589_),
    .B(_09591_),
    .C(_09593_),
    .D(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__nand2_2 _13873_ (.A(\res_h_counter[2] ),
    .B(\res_h_counter[3] ),
    .Y(_09599_));
 sky130_fd_sc_hd__nor2_4 _13874_ (.A(_09561_),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__inv_4 _13875_ (.A(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__nor2_1 _13876_ (.A(_09554_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__inv_2 _13877_ (.A(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__inv_2 _13878_ (.A(_09599_),
    .Y(_09604_));
 sky130_fd_sc_hd__nand2_4 _13879_ (.A(_09556_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__or2_1 _13880_ (.A(_09555_),
    .B(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__nand2_4 _13881_ (.A(_09566_),
    .B(_09604_),
    .Y(_09607_));
 sky130_fd_sc_hd__or2_1 _13882_ (.A(_09555_),
    .B(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__nand2_4 _13883_ (.A(_09604_),
    .B(_09571_),
    .Y(_09609_));
 sky130_fd_sc_hd__or2_1 _13884_ (.A(_09609_),
    .B(_09555_),
    .X(_09610_));
 sky130_fd_sc_hd__clkbuf_8 _13885_ (.A(_09583_),
    .X(_09611_));
 sky130_fd_sc_hd__a41o_1 _13886_ (.A1(_09603_),
    .A2(_09606_),
    .A3(_09608_),
    .A4(_09610_),
    .B1(_09611_),
    .X(_09612_));
 sky130_fd_sc_hd__and4_1 _13887_ (.A(_09574_),
    .B(_09586_),
    .C(_09598_),
    .D(_09612_),
    .X(_09613_));
 sky130_fd_sc_hd__o21ai_1 _13888_ (.A1(_09548_),
    .A2(_09550_),
    .B1(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__a211o_1 _13889_ (.A1(_09533_),
    .A2(_09540_),
    .B1(_09544_),
    .C1(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__buf_8 _13890_ (.A(_08995_),
    .X(_09616_));
 sky130_fd_sc_hd__and3_2 _13891_ (.A(_09542_),
    .B(_09013_),
    .C(_09035_),
    .X(_09617_));
 sky130_fd_sc_hd__clkinv_4 _13892_ (.A(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__or3_1 _13893_ (.A(_09616_),
    .B(_09559_),
    .C(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__inv_2 _13894_ (.A(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__buf_6 _13895_ (.A(_09617_),
    .X(_09621_));
 sky130_fd_sc_hd__and3_1 _13896_ (.A(_09621_),
    .B(_09563_),
    .C(_09551_),
    .X(_09622_));
 sky130_fd_sc_hd__clkbuf_4 _13897_ (.A(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__nor2_2 _13898_ (.A(_09567_),
    .B(_09618_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand2_1 _13899_ (.A(_09624_),
    .B(_09546_),
    .Y(_09625_));
 sky130_fd_sc_hd__nor2_2 _13900_ (.A(_09572_),
    .B(_09618_),
    .Y(_09626_));
 sky130_fd_sc_hd__nand2_1 _13901_ (.A(_09626_),
    .B(_09546_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand2_1 _13902_ (.A(_09625_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__nor2_1 _13903_ (.A(_09588_),
    .B(_09618_),
    .Y(_09629_));
 sky130_fd_sc_hd__nand2_1 _13904_ (.A(_09629_),
    .B(_09546_),
    .Y(_09630_));
 sky130_fd_sc_hd__nor2_4 _13905_ (.A(_09594_),
    .B(_09618_),
    .Y(_09631_));
 sky130_fd_sc_hd__nand2_1 _13906_ (.A(_09631_),
    .B(_09583_),
    .Y(_09632_));
 sky130_fd_sc_hd__nand2_1 _13907_ (.A(_09630_),
    .B(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__clkinv_4 _13908_ (.A(_09590_),
    .Y(_09634_));
 sky130_fd_sc_hd__and3_1 _13909_ (.A(_09621_),
    .B(_09634_),
    .C(_08993_),
    .X(_09635_));
 sky130_fd_sc_hd__clkbuf_4 _13910_ (.A(_09635_),
    .X(_09636_));
 sky130_fd_sc_hd__inv_2 _13911_ (.A(_09592_),
    .Y(_09637_));
 sky130_fd_sc_hd__and3_1 _13912_ (.A(_09621_),
    .B(_09637_),
    .C(_09541_),
    .X(_09638_));
 sky130_fd_sc_hd__clkbuf_4 _13913_ (.A(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__or2_1 _13914_ (.A(_09636_),
    .B(_09639_),
    .X(_09640_));
 sky130_fd_sc_hd__or2_1 _13915_ (.A(_09633_),
    .B(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__or4_1 _13916_ (.A(_09620_),
    .B(_09623_),
    .C(_09628_),
    .D(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__inv_2 _13917_ (.A(_09607_),
    .Y(_09643_));
 sky130_fd_sc_hd__and3_1 _13918_ (.A(_09621_),
    .B(_09545_),
    .C(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__buf_2 _13919_ (.A(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__clkinv_4 _13920_ (.A(_09609_),
    .Y(_09646_));
 sky130_fd_sc_hd__and3_1 _13921_ (.A(_09621_),
    .B(_09646_),
    .C(_09551_),
    .X(_09647_));
 sky130_fd_sc_hd__clkbuf_4 _13922_ (.A(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__nor2_1 _13923_ (.A(_09605_),
    .B(_09618_),
    .Y(_09649_));
 sky130_fd_sc_hd__nand2_2 _13924_ (.A(_09649_),
    .B(_09611_),
    .Y(_09650_));
 sky130_fd_sc_hd__nor2_1 _13925_ (.A(_09601_),
    .B(_09618_),
    .Y(_09651_));
 sky130_fd_sc_hd__nand2_1 _13926_ (.A(_09651_),
    .B(_09611_),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2_1 _13927_ (.A(_09650_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__and3_1 _13928_ (.A(_09621_),
    .B(_09541_),
    .C(_09577_),
    .X(_09654_));
 sky130_fd_sc_hd__clkbuf_4 _13929_ (.A(_09654_),
    .X(_09655_));
 sky130_fd_sc_hd__clkinv_4 _13930_ (.A(_09584_),
    .Y(_09656_));
 sky130_fd_sc_hd__and3_1 _13931_ (.A(_09621_),
    .B(_09656_),
    .C(_09541_),
    .X(_09657_));
 sky130_fd_sc_hd__clkbuf_4 _13932_ (.A(_09657_),
    .X(_09658_));
 sky130_fd_sc_hd__clkinv_4 _13933_ (.A(_09581_),
    .Y(_09659_));
 sky130_fd_sc_hd__and3_1 _13934_ (.A(_09621_),
    .B(_09659_),
    .C(_09541_),
    .X(_09660_));
 sky130_fd_sc_hd__clkbuf_4 _13935_ (.A(_09660_),
    .X(_09661_));
 sky130_fd_sc_hd__clkinv_4 _13936_ (.A(_09579_),
    .Y(_09662_));
 sky130_fd_sc_hd__and3_4 _13937_ (.A(_09621_),
    .B(_09662_),
    .C(_09541_),
    .X(_09663_));
 sky130_fd_sc_hd__or4_1 _13938_ (.A(_09655_),
    .B(_09658_),
    .C(_09661_),
    .D(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__or4_1 _13939_ (.A(_09645_),
    .B(_09648_),
    .C(_09653_),
    .D(_09664_),
    .X(_09665_));
 sky130_fd_sc_hd__nor2_1 _13940_ (.A(_09642_),
    .B(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__and3_1 _13941_ (.A(_09536_),
    .B(_09013_),
    .C(_09035_),
    .X(_09667_));
 sky130_fd_sc_hd__buf_6 _13942_ (.A(_09667_),
    .X(_09668_));
 sky130_fd_sc_hd__nand2_1 _13943_ (.A(_09668_),
    .B(_09541_),
    .Y(_09669_));
 sky130_fd_sc_hd__and3_1 _13944_ (.A(_09553_),
    .B(_09013_),
    .C(_09035_),
    .X(_09670_));
 sky130_fd_sc_hd__buf_6 _13945_ (.A(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__clkbuf_4 _13946_ (.A(_09671_),
    .X(_09672_));
 sky130_fd_sc_hd__clkinv_4 _13947_ (.A(_09572_),
    .Y(_09673_));
 sky130_fd_sc_hd__and3_1 _13948_ (.A(_09672_),
    .B(_09673_),
    .C(_09545_),
    .X(_09674_));
 sky130_fd_sc_hd__clkbuf_4 _13949_ (.A(_09674_),
    .X(_09675_));
 sky130_fd_sc_hd__and3_4 _13950_ (.A(_09672_),
    .B(_09551_),
    .C(_09568_),
    .X(_09676_));
 sky130_fd_sc_hd__and3_4 _13951_ (.A(_09672_),
    .B(_09551_),
    .C(_09558_),
    .X(_09677_));
 sky130_fd_sc_hd__and3_4 _13952_ (.A(_09672_),
    .B(_09563_),
    .C(_09551_),
    .X(_09678_));
 sky130_fd_sc_hd__or2_1 _13953_ (.A(_09677_),
    .B(_09678_),
    .X(_09679_));
 sky130_fd_sc_hd__or3_1 _13954_ (.A(_09675_),
    .B(_09676_),
    .C(_09679_),
    .X(_09680_));
 sky130_fd_sc_hd__clkinv_4 _13955_ (.A(_09588_),
    .Y(_09681_));
 sky130_fd_sc_hd__and3_4 _13956_ (.A(_09672_),
    .B(_09681_),
    .C(_09583_),
    .X(_09682_));
 sky130_fd_sc_hd__inv_4 _13957_ (.A(_09594_),
    .Y(_09683_));
 sky130_fd_sc_hd__and3_1 _13958_ (.A(_09672_),
    .B(_09545_),
    .C(_09683_),
    .X(_09684_));
 sky130_fd_sc_hd__clkbuf_4 _13959_ (.A(_09684_),
    .X(_09685_));
 sky130_fd_sc_hd__inv_2 _13960_ (.A(_09671_),
    .Y(_09686_));
 sky130_fd_sc_hd__nor2_2 _13961_ (.A(_09592_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand2_1 _13962_ (.A(_09687_),
    .B(_09546_),
    .Y(_09688_));
 sky130_fd_sc_hd__inv_2 _13963_ (.A(_09688_),
    .Y(_09689_));
 sky130_fd_sc_hd__nor2_1 _13964_ (.A(_09590_),
    .B(_09686_),
    .Y(_09690_));
 sky130_fd_sc_hd__buf_4 _13965_ (.A(_09583_),
    .X(_09691_));
 sky130_fd_sc_hd__nand2_1 _13966_ (.A(_09690_),
    .B(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__inv_2 _13967_ (.A(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__or4_1 _13968_ (.A(_09682_),
    .B(_09685_),
    .C(_09689_),
    .D(_09693_),
    .X(_09694_));
 sky130_fd_sc_hd__nor2_2 _13969_ (.A(_09601_),
    .B(_09686_),
    .Y(_09695_));
 sky130_fd_sc_hd__and3_1 _13970_ (.A(_09672_),
    .B(_09646_),
    .C(_09541_),
    .X(_09696_));
 sky130_fd_sc_hd__buf_2 _13971_ (.A(_09696_),
    .X(_09697_));
 sky130_fd_sc_hd__and3_1 _13972_ (.A(_09672_),
    .B(_09541_),
    .C(_09643_),
    .X(_09698_));
 sky130_fd_sc_hd__buf_2 _13973_ (.A(_09698_),
    .X(_09699_));
 sky130_fd_sc_hd__nor2_1 _13974_ (.A(_09605_),
    .B(_09686_),
    .Y(_09700_));
 sky130_fd_sc_hd__inv_2 _13975_ (.A(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__nor2_4 _13976_ (.A(_09531_),
    .B(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__a2111o_1 _13977_ (.A1(_09611_),
    .A2(_09695_),
    .B1(_09697_),
    .C1(_09699_),
    .D1(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__and3_1 _13978_ (.A(_09672_),
    .B(_09577_),
    .C(_09545_),
    .X(_09704_));
 sky130_fd_sc_hd__clkbuf_4 _13979_ (.A(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__and3_1 _13980_ (.A(_09672_),
    .B(_09545_),
    .C(_09662_),
    .X(_09706_));
 sky130_fd_sc_hd__clkbuf_4 _13981_ (.A(_09706_),
    .X(_09707_));
 sky130_fd_sc_hd__and3_4 _13982_ (.A(_09672_),
    .B(_09551_),
    .C(_09659_),
    .X(_09708_));
 sky130_fd_sc_hd__and3_4 _13983_ (.A(_09672_),
    .B(_09656_),
    .C(_09551_),
    .X(_09709_));
 sky130_fd_sc_hd__or2_1 _13984_ (.A(_09708_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__nor3_1 _13985_ (.A(_09705_),
    .B(_09707_),
    .C(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__or2b_1 _13986_ (.A(_09703_),
    .B_N(_09711_),
    .X(_09712_));
 sky130_fd_sc_hd__nor3_1 _13987_ (.A(_09680_),
    .B(_09694_),
    .C(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__and3_2 _13988_ (.A(_09549_),
    .B(_09013_),
    .C(_09035_),
    .X(_09714_));
 sky130_fd_sc_hd__buf_4 _13989_ (.A(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__and3_4 _13990_ (.A(_09715_),
    .B(_09583_),
    .C(_09577_),
    .X(_09716_));
 sky130_fd_sc_hd__and3_1 _13991_ (.A(_09715_),
    .B(_09656_),
    .C(_09545_),
    .X(_09717_));
 sky130_fd_sc_hd__clkbuf_4 _13992_ (.A(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__and3_1 _13993_ (.A(_09715_),
    .B(_09659_),
    .C(_09545_),
    .X(_09719_));
 sky130_fd_sc_hd__clkbuf_4 _13994_ (.A(_09719_),
    .X(_09720_));
 sky130_fd_sc_hd__and3_4 _13995_ (.A(_09715_),
    .B(_09662_),
    .C(_09583_),
    .X(_09721_));
 sky130_fd_sc_hd__or4_1 _13996_ (.A(_09716_),
    .B(_09718_),
    .C(_09720_),
    .D(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__inv_2 _13997_ (.A(_09714_),
    .Y(_09723_));
 sky130_fd_sc_hd__nor2_1 _13998_ (.A(_09588_),
    .B(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__and3_1 _13999_ (.A(_09715_),
    .B(_09634_),
    .C(_09545_),
    .X(_09725_));
 sky130_fd_sc_hd__clkbuf_4 _14000_ (.A(_09725_),
    .X(_09726_));
 sky130_fd_sc_hd__and3_1 _14001_ (.A(_09715_),
    .B(_09637_),
    .C(_09545_),
    .X(_09727_));
 sky130_fd_sc_hd__clkbuf_4 _14002_ (.A(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__and3_1 _14003_ (.A(_09715_),
    .B(_09683_),
    .C(_09583_),
    .X(_09729_));
 sky130_fd_sc_hd__clkbuf_4 _14004_ (.A(_09729_),
    .X(_09730_));
 sky130_fd_sc_hd__a2111oi_1 _14005_ (.A1(_09547_),
    .A2(_09724_),
    .B1(_09726_),
    .C1(_09728_),
    .D1(_09730_),
    .Y(_09731_));
 sky130_fd_sc_hd__nor2_1 _14006_ (.A(_09567_),
    .B(_09723_),
    .Y(_09732_));
 sky130_fd_sc_hd__nand2_1 _14007_ (.A(_09732_),
    .B(_09583_),
    .Y(_09733_));
 sky130_fd_sc_hd__nor2_1 _14008_ (.A(_09559_),
    .B(_09723_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_1 _14009_ (.A(_09734_),
    .B(_09691_),
    .Y(_09735_));
 sky130_fd_sc_hd__nor2_1 _14010_ (.A(_09564_),
    .B(_09723_),
    .Y(_09736_));
 sky130_fd_sc_hd__nand2_1 _14011_ (.A(_09736_),
    .B(_09691_),
    .Y(_09737_));
 sky130_fd_sc_hd__nor2_1 _14012_ (.A(_09572_),
    .B(_09723_),
    .Y(_09738_));
 sky130_fd_sc_hd__nand2_1 _14013_ (.A(_09738_),
    .B(_09583_),
    .Y(_09739_));
 sky130_fd_sc_hd__and4_1 _14014_ (.A(_09733_),
    .B(_09735_),
    .C(_09737_),
    .D(_09739_),
    .X(_09740_));
 sky130_fd_sc_hd__nand2_1 _14015_ (.A(_09731_),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__and3_2 _14016_ (.A(_09715_),
    .B(_09646_),
    .C(_09545_),
    .X(_09742_));
 sky130_fd_sc_hd__and3_2 _14017_ (.A(_09715_),
    .B(_09545_),
    .C(_09643_),
    .X(_09743_));
 sky130_fd_sc_hd__nor2_1 _14018_ (.A(_09601_),
    .B(_09723_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_1 _14019_ (.A(_09744_),
    .B(_09546_),
    .Y(_09745_));
 sky130_fd_sc_hd__inv_2 _14020_ (.A(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__or3_4 _14021_ (.A(_09530_),
    .B(_09605_),
    .C(_09723_),
    .X(_09747_));
 sky130_fd_sc_hd__or4b_1 _14022_ (.A(_09742_),
    .B(_09743_),
    .C(_09746_),
    .D_N(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__nor3_1 _14023_ (.A(_09722_),
    .B(_09741_),
    .C(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__and4_1 _14024_ (.A(_09666_),
    .B(_09669_),
    .C(_09713_),
    .D(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__and3_4 _14025_ (.A(_09549_),
    .B(_09013_),
    .C(\res_h_counter[7] ),
    .X(_09751_));
 sky130_fd_sc_hd__inv_12 _14026_ (.A(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__and3_4 _14027_ (.A(_09542_),
    .B(_09013_),
    .C(\res_h_counter[7] ),
    .X(_09753_));
 sky130_fd_sc_hd__inv_12 _14028_ (.A(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__and3_4 _14029_ (.A(_09553_),
    .B(_09013_),
    .C(\res_h_counter[7] ),
    .X(_09755_));
 sky130_fd_sc_hd__inv_12 _14030_ (.A(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__and3_1 _14031_ (.A(_09536_),
    .B(_09013_),
    .C(\res_h_counter[7] ),
    .X(_09757_));
 sky130_fd_sc_hd__buf_4 _14032_ (.A(_09757_),
    .X(_09758_));
 sky130_fd_sc_hd__inv_2 _14033_ (.A(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__clkbuf_16 _14034_ (.A(_09759_),
    .X(_09760_));
 sky130_fd_sc_hd__a41o_1 _14035_ (.A1(_09752_),
    .A2(_09754_),
    .A3(_09756_),
    .A4(_09760_),
    .B1(_09548_),
    .X(_09761_));
 sky130_fd_sc_hd__nor2_8 _14036_ (.A(\res_h_counter[7] ),
    .B(_09013_),
    .Y(_09762_));
 sky130_fd_sc_hd__nand2_4 _14037_ (.A(_09542_),
    .B(_09762_),
    .Y(_09763_));
 sky130_fd_sc_hd__buf_12 _14038_ (.A(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__nand2_8 _14039_ (.A(_09549_),
    .B(_09762_),
    .Y(_09765_));
 sky130_fd_sc_hd__nand2_8 _14040_ (.A(_09762_),
    .B(_09536_),
    .Y(_09766_));
 sky130_fd_sc_hd__nand2_4 _14041_ (.A(_09762_),
    .B(_09553_),
    .Y(_09767_));
 sky130_fd_sc_hd__clkbuf_16 _14042_ (.A(_09767_),
    .X(_09768_));
 sky130_fd_sc_hd__a41o_1 _14043_ (.A1(_09764_),
    .A2(_09765_),
    .A3(_09766_),
    .A4(_09768_),
    .B1(_09548_),
    .X(_09769_));
 sky130_fd_sc_hd__and2_1 _14044_ (.A(_09761_),
    .B(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__nand3b_2 _14045_ (.A_N(_09615_),
    .B(_09750_),
    .C(_09770_),
    .Y(_09771_));
 sky130_fd_sc_hd__and3_1 _14046_ (.A(_09714_),
    .B(_09634_),
    .C(_08995_),
    .X(_09772_));
 sky130_fd_sc_hd__clkbuf_4 _14047_ (.A(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__and3_1 _14048_ (.A(_09715_),
    .B(_09683_),
    .C(_08995_),
    .X(_09774_));
 sky130_fd_sc_hd__buf_4 _14049_ (.A(_09774_),
    .X(_09775_));
 sky130_fd_sc_hd__nand2_2 _14050_ (.A(_09724_),
    .B(_09616_),
    .Y(_09776_));
 sky130_fd_sc_hd__clkinv_4 _14051_ (.A(_09776_),
    .Y(_09777_));
 sky130_fd_sc_hd__clkbuf_8 _14052_ (.A(_08994_),
    .X(_09778_));
 sky130_fd_sc_hd__and3_1 _14053_ (.A(_09715_),
    .B(_09637_),
    .C(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__clkbuf_8 _14054_ (.A(_09779_),
    .X(_09780_));
 sky130_fd_sc_hd__or4_1 _14055_ (.A(_09773_),
    .B(_09775_),
    .C(_09777_),
    .D(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__and3_1 _14056_ (.A(_09714_),
    .B(_08995_),
    .C(_09577_),
    .X(_09782_));
 sky130_fd_sc_hd__buf_4 _14057_ (.A(_09782_),
    .X(_09783_));
 sky130_fd_sc_hd__and3_1 _14058_ (.A(_09715_),
    .B(_09656_),
    .C(_08995_),
    .X(_09784_));
 sky130_fd_sc_hd__clkbuf_8 _14059_ (.A(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__and3_1 _14060_ (.A(_09715_),
    .B(_09662_),
    .C(_09778_),
    .X(_09786_));
 sky130_fd_sc_hd__clkbuf_4 _14061_ (.A(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__and3_1 _14062_ (.A(_09715_),
    .B(_09659_),
    .C(_09778_),
    .X(_09788_));
 sky130_fd_sc_hd__clkbuf_4 _14063_ (.A(_09788_),
    .X(_09789_));
 sky130_fd_sc_hd__or4_1 _14064_ (.A(_09783_),
    .B(_09785_),
    .C(_09787_),
    .D(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__nand2_2 _14065_ (.A(_09738_),
    .B(_09616_),
    .Y(_09791_));
 sky130_fd_sc_hd__clkinv_4 _14066_ (.A(_09791_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_2 _14067_ (.A(_09736_),
    .B(_09616_),
    .Y(_09793_));
 sky130_fd_sc_hd__clkinv_4 _14068_ (.A(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_2 _14069_ (.A(_09732_),
    .B(_09616_),
    .Y(_09795_));
 sky130_fd_sc_hd__clkinv_4 _14070_ (.A(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__nand2_2 _14071_ (.A(_09734_),
    .B(_09616_),
    .Y(_09797_));
 sky130_fd_sc_hd__clkinv_4 _14072_ (.A(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__or4_1 _14073_ (.A(_09792_),
    .B(_09794_),
    .C(_09796_),
    .D(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__and3_1 _14074_ (.A(_09715_),
    .B(_09646_),
    .C(_09778_),
    .X(_09800_));
 sky130_fd_sc_hd__clkbuf_8 _14075_ (.A(_09800_),
    .X(_09801_));
 sky130_fd_sc_hd__and3_1 _14076_ (.A(_09715_),
    .B(_09530_),
    .C(_09643_),
    .X(_09802_));
 sky130_fd_sc_hd__buf_2 _14077_ (.A(_09802_),
    .X(_09803_));
 sky130_fd_sc_hd__nor3_4 _14078_ (.A(_09541_),
    .B(_09605_),
    .C(_09723_),
    .Y(_09804_));
 sky130_fd_sc_hd__nand2_1 _14079_ (.A(_09744_),
    .B(_09531_),
    .Y(_09805_));
 sky130_fd_sc_hd__inv_2 _14080_ (.A(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__or4_1 _14081_ (.A(_09801_),
    .B(_09803_),
    .C(_09804_),
    .D(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__or4_1 _14082_ (.A(_09781_),
    .B(_09790_),
    .C(_09799_),
    .D(_09807_),
    .X(_09808_));
 sky130_fd_sc_hd__and3_4 _14083_ (.A(_09671_),
    .B(_09681_),
    .C(_09530_),
    .X(_09809_));
 sky130_fd_sc_hd__and3_1 _14084_ (.A(_09671_),
    .B(_09778_),
    .C(_09683_),
    .X(_09810_));
 sky130_fd_sc_hd__buf_6 _14085_ (.A(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__nand2_2 _14086_ (.A(_09690_),
    .B(_09616_),
    .Y(_09812_));
 sky130_fd_sc_hd__inv_2 _14087_ (.A(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_1 _14088_ (.A(_09687_),
    .B(_09616_),
    .Y(_09814_));
 sky130_fd_sc_hd__inv_2 _14089_ (.A(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__or4_1 _14090_ (.A(_09809_),
    .B(_09811_),
    .C(_09813_),
    .D(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__and3_2 _14091_ (.A(_09671_),
    .B(_09646_),
    .C(_09530_),
    .X(_09817_));
 sky130_fd_sc_hd__and3_1 _14092_ (.A(_09671_),
    .B(_09778_),
    .C(_09643_),
    .X(_09818_));
 sky130_fd_sc_hd__buf_2 _14093_ (.A(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__nand2_1 _14094_ (.A(_09695_),
    .B(_09530_),
    .Y(_09820_));
 sky130_fd_sc_hd__inv_2 _14095_ (.A(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__nor2_4 _14096_ (.A(_09545_),
    .B(_09701_),
    .Y(_09822_));
 sky130_fd_sc_hd__or4_1 _14097_ (.A(_09817_),
    .B(_09819_),
    .C(_09821_),
    .D(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__and3_4 _14098_ (.A(_09671_),
    .B(_09673_),
    .C(_09530_),
    .X(_09824_));
 sky130_fd_sc_hd__and3_1 _14099_ (.A(_09671_),
    .B(_09778_),
    .C(_09568_),
    .X(_09825_));
 sky130_fd_sc_hd__clkbuf_4 _14100_ (.A(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__and3_4 _14101_ (.A(_09671_),
    .B(_09616_),
    .C(_09558_),
    .X(_09827_));
 sky130_fd_sc_hd__and3_4 _14102_ (.A(_09672_),
    .B(_09563_),
    .C(_09616_),
    .X(_09828_));
 sky130_fd_sc_hd__or4_1 _14103_ (.A(_09824_),
    .B(_09826_),
    .C(_09827_),
    .D(_09828_),
    .X(_09829_));
 sky130_fd_sc_hd__and3_2 _14104_ (.A(_09672_),
    .B(_09577_),
    .C(_09616_),
    .X(_09830_));
 sky130_fd_sc_hd__and3_1 _14105_ (.A(_09671_),
    .B(_09530_),
    .C(_09659_),
    .X(_09831_));
 sky130_fd_sc_hd__buf_2 _14106_ (.A(_09831_),
    .X(_09832_));
 sky130_fd_sc_hd__and3_2 _14107_ (.A(_09672_),
    .B(_09656_),
    .C(_09616_),
    .X(_09833_));
 sky130_fd_sc_hd__and3_2 _14108_ (.A(_09672_),
    .B(_09616_),
    .C(_09662_),
    .X(_09834_));
 sky130_fd_sc_hd__or4_1 _14109_ (.A(_09830_),
    .B(_09832_),
    .C(_09833_),
    .D(_09834_),
    .X(_09835_));
 sky130_fd_sc_hd__or4_1 _14110_ (.A(_09816_),
    .B(_09823_),
    .C(_09829_),
    .D(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__inv_6 _14111_ (.A(_09668_),
    .Y(_09837_));
 sky130_fd_sc_hd__nor2_1 _14112_ (.A(_09559_),
    .B(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__nor2_1 _14113_ (.A(_09567_),
    .B(_09837_),
    .Y(_09839_));
 sky130_fd_sc_hd__nor2_4 _14114_ (.A(_09564_),
    .B(_09837_),
    .Y(_09840_));
 sky130_fd_sc_hd__o31a_1 _14115_ (.A1(_09838_),
    .A2(_09839_),
    .A3(_09840_),
    .B1(_09531_),
    .X(_09841_));
 sky130_fd_sc_hd__and3_2 _14116_ (.A(_09668_),
    .B(_09634_),
    .C(_08995_),
    .X(_09842_));
 sky130_fd_sc_hd__and3_1 _14117_ (.A(_09668_),
    .B(_08994_),
    .C(_09683_),
    .X(_09843_));
 sky130_fd_sc_hd__buf_6 _14118_ (.A(_09843_),
    .X(_09844_));
 sky130_fd_sc_hd__nor2_1 _14119_ (.A(_09592_),
    .B(_09837_),
    .Y(_09845_));
 sky130_fd_sc_hd__nand2_1 _14120_ (.A(_09845_),
    .B(_09778_),
    .Y(_09846_));
 sky130_fd_sc_hd__inv_2 _14121_ (.A(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__nor2_4 _14122_ (.A(_09588_),
    .B(_09837_),
    .Y(_09848_));
 sky130_fd_sc_hd__nand2_1 _14123_ (.A(_09848_),
    .B(_09530_),
    .Y(_09849_));
 sky130_fd_sc_hd__inv_2 _14124_ (.A(_09849_),
    .Y(_09850_));
 sky130_fd_sc_hd__or4_1 _14125_ (.A(_09842_),
    .B(_09844_),
    .C(_09847_),
    .D(_09850_),
    .X(_09851_));
 sky130_fd_sc_hd__and3_1 _14126_ (.A(_09668_),
    .B(_09659_),
    .C(_08994_),
    .X(_09852_));
 sky130_fd_sc_hd__clkbuf_4 _14127_ (.A(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__and3_1 _14128_ (.A(_09668_),
    .B(_09577_),
    .C(_08994_),
    .X(_09854_));
 sky130_fd_sc_hd__clkbuf_4 _14129_ (.A(_09854_),
    .X(_09855_));
 sky130_fd_sc_hd__and3_1 _14130_ (.A(_09668_),
    .B(_08994_),
    .C(_09662_),
    .X(_09856_));
 sky130_fd_sc_hd__clkbuf_4 _14131_ (.A(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__nor2_4 _14132_ (.A(_09584_),
    .B(_09837_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand2_1 _14133_ (.A(_09858_),
    .B(_09778_),
    .Y(_09859_));
 sky130_fd_sc_hd__inv_2 _14134_ (.A(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__or4_1 _14135_ (.A(_09853_),
    .B(_09855_),
    .C(_09857_),
    .D(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__nor2_4 _14136_ (.A(_09609_),
    .B(_09837_),
    .Y(_09862_));
 sky130_fd_sc_hd__nand2_1 _14137_ (.A(_09862_),
    .B(_09778_),
    .Y(_09863_));
 sky130_fd_sc_hd__inv_2 _14138_ (.A(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__nor2_1 _14139_ (.A(_09601_),
    .B(_09837_),
    .Y(_09865_));
 sky130_fd_sc_hd__nand2_1 _14140_ (.A(_09865_),
    .B(_09530_),
    .Y(_09866_));
 sky130_fd_sc_hd__inv_2 _14141_ (.A(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__nor2_1 _14142_ (.A(_09605_),
    .B(_09837_),
    .Y(_09868_));
 sky130_fd_sc_hd__nand2_1 _14143_ (.A(_09868_),
    .B(_09530_),
    .Y(_09869_));
 sky130_fd_sc_hd__inv_4 _14144_ (.A(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__nor2_2 _14145_ (.A(_09607_),
    .B(_09837_),
    .Y(_09871_));
 sky130_fd_sc_hd__nand2_1 _14146_ (.A(_09871_),
    .B(_09778_),
    .Y(_09872_));
 sky130_fd_sc_hd__inv_4 _14147_ (.A(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__or4_1 _14148_ (.A(_09864_),
    .B(_09867_),
    .C(_09870_),
    .D(_09873_),
    .X(_09874_));
 sky130_fd_sc_hd__or4_1 _14149_ (.A(_09841_),
    .B(_09851_),
    .C(_09861_),
    .D(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__and3_1 _14150_ (.A(_09621_),
    .B(_09563_),
    .C(_08995_),
    .X(_09876_));
 sky130_fd_sc_hd__clkbuf_4 _14151_ (.A(_09876_),
    .X(_09877_));
 sky130_fd_sc_hd__and3_4 _14152_ (.A(_09621_),
    .B(_09558_),
    .C(_09778_),
    .X(_09878_));
 sky130_fd_sc_hd__nand2_1 _14153_ (.A(_09624_),
    .B(_09616_),
    .Y(_09879_));
 sky130_fd_sc_hd__nand2_1 _14154_ (.A(_09626_),
    .B(_09616_),
    .Y(_09880_));
 sky130_fd_sc_hd__nand2_1 _14155_ (.A(_09879_),
    .B(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__or3_1 _14156_ (.A(_09877_),
    .B(_09878_),
    .C(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__and3_1 _14157_ (.A(_09621_),
    .B(_09637_),
    .C(_08995_),
    .X(_09883_));
 sky130_fd_sc_hd__clkbuf_4 _14158_ (.A(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__and3_1 _14159_ (.A(_09621_),
    .B(_09634_),
    .C(_08995_),
    .X(_09885_));
 sky130_fd_sc_hd__clkbuf_4 _14160_ (.A(_09885_),
    .X(_09886_));
 sky130_fd_sc_hd__and3_1 _14161_ (.A(_09621_),
    .B(_09778_),
    .C(_09681_),
    .X(_09887_));
 sky130_fd_sc_hd__buf_2 _14162_ (.A(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__a2111o_1 _14163_ (.A1(_09531_),
    .A2(_09631_),
    .B1(_09884_),
    .C1(_09886_),
    .D1(_09888_),
    .X(_09889_));
 sky130_fd_sc_hd__and3_4 _14164_ (.A(_09621_),
    .B(_09656_),
    .C(_08995_),
    .X(_09890_));
 sky130_fd_sc_hd__and3_1 _14165_ (.A(_09617_),
    .B(_09662_),
    .C(_08994_),
    .X(_09891_));
 sky130_fd_sc_hd__buf_4 _14166_ (.A(_09891_),
    .X(_09892_));
 sky130_fd_sc_hd__nor2_1 _14167_ (.A(_09576_),
    .B(_09618_),
    .Y(_09893_));
 sky130_fd_sc_hd__nand2_1 _14168_ (.A(_09893_),
    .B(_09778_),
    .Y(_09894_));
 sky130_fd_sc_hd__inv_4 _14169_ (.A(_09894_),
    .Y(_09895_));
 sky130_fd_sc_hd__and3_4 _14170_ (.A(_09621_),
    .B(_09659_),
    .C(_09778_),
    .X(_09896_));
 sky130_fd_sc_hd__or4_1 _14171_ (.A(_09890_),
    .B(_09892_),
    .C(_09895_),
    .D(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__nor2_1 _14172_ (.A(_09609_),
    .B(_09618_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand2_1 _14173_ (.A(_09898_),
    .B(_09530_),
    .Y(_09899_));
 sky130_fd_sc_hd__clkinv_4 _14174_ (.A(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__nor2_1 _14175_ (.A(_09607_),
    .B(_09618_),
    .Y(_09901_));
 sky130_fd_sc_hd__nand2_1 _14176_ (.A(_09901_),
    .B(_09530_),
    .Y(_09902_));
 sky130_fd_sc_hd__clkinv_4 _14177_ (.A(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__nand2_1 _14178_ (.A(_09649_),
    .B(_09530_),
    .Y(_09904_));
 sky130_fd_sc_hd__clkinv_4 _14179_ (.A(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand2_1 _14180_ (.A(_09651_),
    .B(_09530_),
    .Y(_09906_));
 sky130_fd_sc_hd__inv_2 _14181_ (.A(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__or4_1 _14182_ (.A(_09900_),
    .B(_09903_),
    .C(_09905_),
    .D(_09907_),
    .X(_09908_));
 sky130_fd_sc_hd__or4_1 _14183_ (.A(_09882_),
    .B(_09889_),
    .C(_09897_),
    .D(_09908_),
    .X(_09909_));
 sky130_fd_sc_hd__or2_1 _14184_ (.A(_09875_),
    .B(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__or3_1 _14185_ (.A(_09808_),
    .B(_09836_),
    .C(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__nor2_2 _14186_ (.A(_09771_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__nand2_1 _14187_ (.A(_09840_),
    .B(_09531_),
    .Y(_09913_));
 sky130_fd_sc_hd__inv_2 _14188_ (.A(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__a22o_1 _14189_ (.A1(_09842_),
    .A2(\line_cache[6][0] ),
    .B1(\line_cache[5][0] ),
    .B2(_09844_),
    .X(_09915_));
 sky130_fd_sc_hd__a221o_1 _14190_ (.A1(\line_cache[4][0] ),
    .A2(_09850_),
    .B1(\line_cache[3][0] ),
    .B2(_09914_),
    .C1(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__buf_4 _14191_ (.A(_09838_),
    .X(_09917_));
 sky130_fd_sc_hd__and3_1 _14192_ (.A(_09917_),
    .B(_09533_),
    .C(\line_cache[2][0] ),
    .X(_09918_));
 sky130_fd_sc_hd__buf_4 _14193_ (.A(_09839_),
    .X(_09919_));
 sky130_fd_sc_hd__and3_1 _14194_ (.A(_09919_),
    .B(_09533_),
    .C(\line_cache[1][0] ),
    .X(_09920_));
 sky130_fd_sc_hd__a211o_1 _14195_ (.A1(\line_cache[15][0] ),
    .A2(_09867_),
    .B1(_09918_),
    .C1(_09920_),
    .X(_09921_));
 sky130_fd_sc_hd__clkbuf_4 _14196_ (.A(_09695_),
    .X(_09922_));
 sky130_fd_sc_hd__and3_1 _14197_ (.A(_09922_),
    .B(_09532_),
    .C(\line_cache[63][0] ),
    .X(_09923_));
 sky130_fd_sc_hd__a31o_1 _14198_ (.A1(_09548_),
    .A2(\line_cache[319][0] ),
    .A3(_09922_),
    .B1(_09923_),
    .X(_09924_));
 sky130_fd_sc_hd__a221o_1 _14199_ (.A1(\line_cache[47][0] ),
    .A2(_09806_),
    .B1(\line_cache[31][0] ),
    .B2(_09907_),
    .C1(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__nor2_4 _14200_ (.A(_09547_),
    .B(_09603_),
    .Y(_09926_));
 sky130_fd_sc_hd__clkinv_4 _14201_ (.A(_09652_),
    .Y(_09927_));
 sky130_fd_sc_hd__nand2_1 _14202_ (.A(_09746_),
    .B(\line_cache[303][0] ),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_1 _14203_ (.A(_09865_),
    .B(_09547_),
    .Y(_09929_));
 sky130_fd_sc_hd__inv_2 _14204_ (.A(_09929_),
    .Y(_09930_));
 sky130_fd_sc_hd__nand2_1 _14205_ (.A(_09930_),
    .B(\line_cache[271][0] ),
    .Y(_09931_));
 sky130_fd_sc_hd__nand2_1 _14206_ (.A(_09928_),
    .B(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__a221oi_2 _14207_ (.A1(\line_cache[255][0] ),
    .A2(_09926_),
    .B1(\line_cache[287][0] ),
    .B2(_09927_),
    .C1(_09932_),
    .Y(_09933_));
 sky130_fd_sc_hd__or4b_1 _14208_ (.A(_09916_),
    .B(_09921_),
    .C(_09925_),
    .D_N(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__a22o_1 _14209_ (.A1(_09803_),
    .A2(\line_cache[45][0] ),
    .B1(\line_cache[46][0] ),
    .B2(_09804_),
    .X(_09935_));
 sky130_fd_sc_hd__a22o_1 _14210_ (.A1(_09824_),
    .A2(\line_cache[48][0] ),
    .B1(\line_cache[49][0] ),
    .B2(_09826_),
    .X(_09936_));
 sky130_fd_sc_hd__nand2_1 _14211_ (.A(_09787_),
    .B(\line_cache[41][0] ),
    .Y(_09937_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(_09789_),
    .B(\line_cache[42][0] ),
    .Y(_09938_));
 sky130_fd_sc_hd__nand2_1 _14213_ (.A(_09937_),
    .B(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__a221oi_4 _14214_ (.A1(_09785_),
    .A2(\line_cache[43][0] ),
    .B1(\line_cache[44][0] ),
    .B2(_09801_),
    .C1(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__or3b_1 _14215_ (.A(_09935_),
    .B(_09936_),
    .C_N(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__a22o_1 _14216_ (.A1(_09699_),
    .A2(\line_cache[317][0] ),
    .B1(\line_cache[316][0] ),
    .B2(_09697_),
    .X(_09942_));
 sky130_fd_sc_hd__a22o_1 _14217_ (.A1(_09832_),
    .A2(\line_cache[58][0] ),
    .B1(\line_cache[59][0] ),
    .B2(_09833_),
    .X(_09943_));
 sky130_fd_sc_hd__a22o_1 _14218_ (.A1(_09819_),
    .A2(\line_cache[61][0] ),
    .B1(\line_cache[60][0] ),
    .B2(_09817_),
    .X(_09944_));
 sky130_fd_sc_hd__a22o_1 _14219_ (.A1(_09822_),
    .A2(\line_cache[62][0] ),
    .B1(\line_cache[318][0] ),
    .B2(_09702_),
    .X(_09945_));
 sky130_fd_sc_hd__or4_1 _14220_ (.A(_09942_),
    .B(_09943_),
    .C(_09944_),
    .D(_09945_),
    .X(_09946_));
 sky130_fd_sc_hd__a22o_1 _14221_ (.A1(_09675_),
    .A2(\line_cache[304][0] ),
    .B1(\line_cache[305][0] ),
    .B2(_09676_),
    .X(_09947_));
 sky130_fd_sc_hd__a22o_1 _14222_ (.A1(_09705_),
    .A2(\line_cache[312][0] ),
    .B1(\line_cache[313][0] ),
    .B2(_09707_),
    .X(_09948_));
 sky130_fd_sc_hd__a22o_1 _14223_ (.A1(_09708_),
    .A2(\line_cache[314][0] ),
    .B1(\line_cache[315][0] ),
    .B2(_09709_),
    .X(_09949_));
 sky130_fd_sc_hd__a22o_1 _14224_ (.A1(_09677_),
    .A2(\line_cache[306][0] ),
    .B1(\line_cache[307][0] ),
    .B2(_09678_),
    .X(_09950_));
 sky130_fd_sc_hd__or4_1 _14225_ (.A(_09947_),
    .B(_09948_),
    .C(_09949_),
    .D(_09950_),
    .X(_09951_));
 sky130_fd_sc_hd__a22o_1 _14226_ (.A1(_09830_),
    .A2(\line_cache[56][0] ),
    .B1(\line_cache[57][0] ),
    .B2(_09834_),
    .X(_09952_));
 sky130_fd_sc_hd__a22o_1 _14227_ (.A1(_09809_),
    .A2(\line_cache[52][0] ),
    .B1(\line_cache[53][0] ),
    .B2(_09811_),
    .X(_09953_));
 sky130_fd_sc_hd__a22o_1 _14228_ (.A1(_09827_),
    .A2(\line_cache[50][0] ),
    .B1(\line_cache[51][0] ),
    .B2(_09828_),
    .X(_09954_));
 sky130_fd_sc_hd__a22o_1 _14229_ (.A1(_09813_),
    .A2(\line_cache[54][0] ),
    .B1(\line_cache[55][0] ),
    .B2(_09815_),
    .X(_09955_));
 sky130_fd_sc_hd__or4_1 _14230_ (.A(_09952_),
    .B(_09953_),
    .C(_09954_),
    .D(_09955_),
    .X(_09956_));
 sky130_fd_sc_hd__or4_2 _14231_ (.A(_09941_),
    .B(_09946_),
    .C(_09951_),
    .D(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__nand2_1 _14232_ (.A(_09864_),
    .B(\line_cache[12][0] ),
    .Y(_09958_));
 sky130_fd_sc_hd__nand2_1 _14233_ (.A(_09860_),
    .B(\line_cache[11][0] ),
    .Y(_09959_));
 sky130_fd_sc_hd__nand2_1 _14234_ (.A(_09958_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__a221oi_2 _14235_ (.A1(_09870_),
    .A2(\line_cache[14][0] ),
    .B1(\line_cache[13][0] ),
    .B2(_09873_),
    .C1(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__nand2_1 _14236_ (.A(_09853_),
    .B(\line_cache[10][0] ),
    .Y(_09962_));
 sky130_fd_sc_hd__nand2_1 _14237_ (.A(_09857_),
    .B(\line_cache[9][0] ),
    .Y(_09963_));
 sky130_fd_sc_hd__nand2_1 _14238_ (.A(_09962_),
    .B(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__a221oi_1 _14239_ (.A1(_09855_),
    .A2(\line_cache[8][0] ),
    .B1(_09847_),
    .B2(\line_cache[7][0] ),
    .C1(_09964_),
    .Y(_09965_));
 sky130_fd_sc_hd__nand2_1 _14240_ (.A(_09961_),
    .B(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__and3_1 _14241_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][0] ),
    .X(_09967_));
 sky130_fd_sc_hd__a22o_1 _14242_ (.A1(_09884_),
    .A2(\line_cache[23][0] ),
    .B1(\line_cache[22][0] ),
    .B2(_09886_),
    .X(_09968_));
 sky130_fd_sc_hd__inv_2 _14243_ (.A(_09879_),
    .Y(_09969_));
 sky130_fd_sc_hd__inv_2 _14244_ (.A(_09880_),
    .Y(_09970_));
 sky130_fd_sc_hd__a22o_1 _14245_ (.A1(_09877_),
    .A2(\line_cache[19][0] ),
    .B1(\line_cache[18][0] ),
    .B2(_09878_),
    .X(_09971_));
 sky130_fd_sc_hd__a221o_1 _14246_ (.A1(\line_cache[17][0] ),
    .A2(_09969_),
    .B1(\line_cache[16][0] ),
    .B2(_09970_),
    .C1(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__a2111o_1 _14247_ (.A1(\line_cache[20][0] ),
    .A2(_09888_),
    .B1(_09967_),
    .C1(_09968_),
    .D1(_09972_),
    .X(_09973_));
 sky130_fd_sc_hd__a22o_1 _14248_ (.A1(_09796_),
    .A2(\line_cache[33][0] ),
    .B1(\line_cache[34][0] ),
    .B2(_09798_),
    .X(_09974_));
 sky130_fd_sc_hd__a221o_1 _14249_ (.A1(\line_cache[36][0] ),
    .A2(_09777_),
    .B1(\line_cache[35][0] ),
    .B2(_09794_),
    .C1(_09974_),
    .X(_09975_));
 sky130_fd_sc_hd__a22o_1 _14250_ (.A1(_09890_),
    .A2(\line_cache[27][0] ),
    .B1(\line_cache[26][0] ),
    .B2(_09896_),
    .X(_09976_));
 sky130_fd_sc_hd__a221oi_1 _14251_ (.A1(\line_cache[25][0] ),
    .A2(_09892_),
    .B1(\line_cache[24][0] ),
    .B2(_09895_),
    .C1(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__a22o_1 _14252_ (.A1(_09903_),
    .A2(\line_cache[29][0] ),
    .B1(\line_cache[28][0] ),
    .B2(_09900_),
    .X(_09978_));
 sky130_fd_sc_hd__a221oi_1 _14253_ (.A1(\line_cache[32][0] ),
    .A2(_09792_),
    .B1(\line_cache[30][0] ),
    .B2(_09905_),
    .C1(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__nand2_1 _14254_ (.A(_09773_),
    .B(\line_cache[38][0] ),
    .Y(_09980_));
 sky130_fd_sc_hd__nand2_1 _14255_ (.A(_09775_),
    .B(\line_cache[37][0] ),
    .Y(_09981_));
 sky130_fd_sc_hd__nand2_1 _14256_ (.A(_09980_),
    .B(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__a221oi_2 _14257_ (.A1(_09783_),
    .A2(\line_cache[40][0] ),
    .B1(\line_cache[39][0] ),
    .B2(_09780_),
    .C1(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__and4b_1 _14258_ (.A_N(_09975_),
    .B(_09977_),
    .C(_09979_),
    .D(_09983_),
    .X(_09984_));
 sky130_fd_sc_hd__or3b_1 _14259_ (.A(_09966_),
    .B(_09973_),
    .C_N(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__nor3_1 _14260_ (.A(_09934_),
    .B(_09957_),
    .C(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__or2_2 _14261_ (.A(_09572_),
    .B(_09669_),
    .X(_09987_));
 sky130_fd_sc_hd__and2b_1 _14262_ (.A_N(_09987_),
    .B(\line_cache[256][0] ),
    .X(_09988_));
 sky130_fd_sc_hd__and2b_1 _14263_ (.A_N(_09747_),
    .B(\line_cache[302][0] ),
    .X(_09989_));
 sky130_fd_sc_hd__a22o_1 _14264_ (.A1(_09742_),
    .A2(\line_cache[300][0] ),
    .B1(\line_cache[301][0] ),
    .B2(_09743_),
    .X(_09990_));
 sky130_fd_sc_hd__or3_1 _14265_ (.A(_09988_),
    .B(_09989_),
    .C(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__and3_1 _14266_ (.A(_09917_),
    .B(_09546_),
    .C(\line_cache[258][0] ),
    .X(_09992_));
 sky130_fd_sc_hd__and3_1 _14267_ (.A(_09848_),
    .B(_09546_),
    .C(\line_cache[260][0] ),
    .X(_09993_));
 sky130_fd_sc_hd__and3_1 _14268_ (.A(_09919_),
    .B(_09546_),
    .C(\line_cache[257][0] ),
    .X(_09994_));
 sky130_fd_sc_hd__and3_1 _14269_ (.A(_09840_),
    .B(_09691_),
    .C(\line_cache[259][0] ),
    .X(_09995_));
 sky130_fd_sc_hd__or4_1 _14270_ (.A(_09992_),
    .B(_09993_),
    .C(_09994_),
    .D(_09995_),
    .X(_09996_));
 sky130_fd_sc_hd__and3_1 _14271_ (.A(_09858_),
    .B(_09611_),
    .C(\line_cache[267][0] ),
    .X(_09997_));
 sky130_fd_sc_hd__and3_2 _14272_ (.A(_09668_),
    .B(_09583_),
    .C(_09662_),
    .X(_09998_));
 sky130_fd_sc_hd__and3_2 _14273_ (.A(_09668_),
    .B(_09659_),
    .C(_09583_),
    .X(_09999_));
 sky130_fd_sc_hd__a22o_1 _14274_ (.A1(_09998_),
    .A2(\line_cache[265][0] ),
    .B1(\line_cache[266][0] ),
    .B2(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__a311o_1 _14275_ (.A1(_09548_),
    .A2(\line_cache[268][0] ),
    .A3(_09862_),
    .B1(_09997_),
    .C1(_10000_),
    .X(_10001_));
 sky130_fd_sc_hd__and3_1 _14276_ (.A(_09668_),
    .B(_09577_),
    .C(_09546_),
    .X(_10002_));
 sky130_fd_sc_hd__buf_2 _14277_ (.A(_10002_),
    .X(_10003_));
 sky130_fd_sc_hd__nand2_1 _14278_ (.A(_09845_),
    .B(_09547_),
    .Y(_10004_));
 sky130_fd_sc_hd__inv_2 _14279_ (.A(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__and3_1 _14280_ (.A(_09668_),
    .B(_09634_),
    .C(_09583_),
    .X(_10006_));
 sky130_fd_sc_hd__buf_2 _14281_ (.A(_10006_),
    .X(_10007_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(_10007_),
    .B(\line_cache[262][0] ),
    .Y(_10008_));
 sky130_fd_sc_hd__and3_1 _14283_ (.A(_09668_),
    .B(_09583_),
    .C(_09683_),
    .X(_10009_));
 sky130_fd_sc_hd__buf_2 _14284_ (.A(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__nand2_1 _14285_ (.A(_10010_),
    .B(\line_cache[261][0] ),
    .Y(_10011_));
 sky130_fd_sc_hd__nand2_1 _14286_ (.A(_10008_),
    .B(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__a221oi_1 _14287_ (.A1(_10003_),
    .A2(\line_cache[264][0] ),
    .B1(_10005_),
    .B2(\line_cache[263][0] ),
    .C1(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__or4b_1 _14288_ (.A(_09991_),
    .B(_09996_),
    .C(_10001_),
    .D_N(_10013_),
    .X(_10014_));
 sky130_fd_sc_hd__a22o_1 _14289_ (.A1(_09682_),
    .A2(\line_cache[308][0] ),
    .B1(\line_cache[309][0] ),
    .B2(_09685_),
    .X(_10015_));
 sky130_fd_sc_hd__a221o_1 _14290_ (.A1(\line_cache[311][0] ),
    .A2(_09689_),
    .B1(\line_cache[310][0] ),
    .B2(_09693_),
    .C1(_10015_),
    .X(_10016_));
 sky130_fd_sc_hd__nand2_1 _14291_ (.A(_09724_),
    .B(_09546_),
    .Y(_10017_));
 sky130_fd_sc_hd__inv_2 _14292_ (.A(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__a22o_1 _14293_ (.A1(_09728_),
    .A2(\line_cache[295][0] ),
    .B1(\line_cache[294][0] ),
    .B2(_09726_),
    .X(_10019_));
 sky130_fd_sc_hd__a221o_1 _14294_ (.A1(\line_cache[293][0] ),
    .A2(_09730_),
    .B1(\line_cache[292][0] ),
    .B2(_10018_),
    .C1(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__a22o_1 _14295_ (.A1(_09716_),
    .A2(\line_cache[296][0] ),
    .B1(\line_cache[297][0] ),
    .B2(_09721_),
    .X(_10021_));
 sky130_fd_sc_hd__a221o_1 _14296_ (.A1(\line_cache[299][0] ),
    .A2(_09718_),
    .B1(\line_cache[298][0] ),
    .B2(_09720_),
    .C1(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__inv_2 _14297_ (.A(_09737_),
    .Y(_10023_));
 sky130_fd_sc_hd__inv_2 _14298_ (.A(_09735_),
    .Y(_10024_));
 sky130_fd_sc_hd__inv_2 _14299_ (.A(_09739_),
    .Y(_10025_));
 sky130_fd_sc_hd__inv_2 _14300_ (.A(_09733_),
    .Y(_10026_));
 sky130_fd_sc_hd__a22o_1 _14301_ (.A1(_10025_),
    .A2(\line_cache[288][0] ),
    .B1(\line_cache[289][0] ),
    .B2(_10026_),
    .X(_10027_));
 sky130_fd_sc_hd__a221o_1 _14302_ (.A1(\line_cache[291][0] ),
    .A2(_10023_),
    .B1(\line_cache[290][0] ),
    .B2(_10024_),
    .C1(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__or4_2 _14303_ (.A(_10016_),
    .B(_10020_),
    .C(_10022_),
    .D(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__nor2_1 _14304_ (.A(_10014_),
    .B(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__nor2_8 _14305_ (.A(_08993_),
    .B(_09607_),
    .Y(_10031_));
 sky130_fd_sc_hd__inv_12 _14306_ (.A(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__nor2_2 _14307_ (.A(_09537_),
    .B(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__nor2_4 _14308_ (.A(_08993_),
    .B(_09584_),
    .Y(_10034_));
 sky130_fd_sc_hd__buf_6 _14309_ (.A(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__and3_1 _14310_ (.A(_10035_),
    .B(\line_cache[203][0] ),
    .C(_09539_),
    .X(_10036_));
 sky130_fd_sc_hd__nor2_4 _14311_ (.A(_09541_),
    .B(_09605_),
    .Y(_10037_));
 sky130_fd_sc_hd__clkbuf_8 _14312_ (.A(_10037_),
    .X(_10038_));
 sky130_fd_sc_hd__and3_1 _14313_ (.A(_10038_),
    .B(\line_cache[206][0] ),
    .C(_09539_),
    .X(_10039_));
 sky130_fd_sc_hd__nand2_8 _14314_ (.A(_09646_),
    .B(_09530_),
    .Y(_10040_));
 sky130_fd_sc_hd__inv_6 _14315_ (.A(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__and3_1 _14316_ (.A(_10041_),
    .B(\line_cache[204][0] ),
    .C(_09539_),
    .X(_10042_));
 sky130_fd_sc_hd__a2111o_1 _14317_ (.A1(\line_cache[205][0] ),
    .A2(_10033_),
    .B1(_10036_),
    .C1(_10039_),
    .D1(_10042_),
    .X(_10043_));
 sky130_fd_sc_hd__nor2_8 _14318_ (.A(_08993_),
    .B(_09590_),
    .Y(_10044_));
 sky130_fd_sc_hd__inv_12 _14319_ (.A(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__nor2_2 _14320_ (.A(_09537_),
    .B(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__nor2_2 _14321_ (.A(_09537_),
    .B(_09596_),
    .Y(_10047_));
 sky130_fd_sc_hd__nand2_8 _14322_ (.A(_09563_),
    .B(_08994_),
    .Y(_10048_));
 sky130_fd_sc_hd__nor2_2 _14323_ (.A(_09537_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_8 _14324_ (.A(_09681_),
    .B(_08995_),
    .Y(_10050_));
 sky130_fd_sc_hd__nor2_2 _14325_ (.A(_09537_),
    .B(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__a22o_1 _14326_ (.A1(_10049_),
    .A2(\line_cache[195][0] ),
    .B1(\line_cache[196][0] ),
    .B2(_10051_),
    .X(_10052_));
 sky130_fd_sc_hd__a221o_1 _14327_ (.A1(\line_cache[198][0] ),
    .A2(_10046_),
    .B1(\line_cache[197][0] ),
    .B2(_10047_),
    .C1(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__nor2_8 _14328_ (.A(_09541_),
    .B(_09581_),
    .Y(_10054_));
 sky130_fd_sc_hd__clkinv_16 _14329_ (.A(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__nor2_2 _14330_ (.A(_09537_),
    .B(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__nor2_4 _14331_ (.A(_09541_),
    .B(_09579_),
    .Y(_10057_));
 sky130_fd_sc_hd__inv_12 _14332_ (.A(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__nor2_2 _14333_ (.A(_09537_),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__nor2_2 _14334_ (.A(_09537_),
    .B(_09578_),
    .Y(_10060_));
 sky130_fd_sc_hd__nor2_8 _14335_ (.A(_08993_),
    .B(_09592_),
    .Y(_10061_));
 sky130_fd_sc_hd__clkinv_16 _14336_ (.A(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__nor2_2 _14337_ (.A(_09537_),
    .B(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__a22o_1 _14338_ (.A1(_10060_),
    .A2(\line_cache[200][0] ),
    .B1(_10063_),
    .B2(\line_cache[199][0] ),
    .X(_10064_));
 sky130_fd_sc_hd__a221o_1 _14339_ (.A1(\line_cache[202][0] ),
    .A2(_10056_),
    .B1(\line_cache[201][0] ),
    .B2(_10059_),
    .C1(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__inv_2 _14340_ (.A(_09650_),
    .Y(_10066_));
 sky130_fd_sc_hd__inv_4 _14341_ (.A(_09569_),
    .Y(_10067_));
 sky130_fd_sc_hd__and3_1 _14342_ (.A(_10067_),
    .B(\line_cache[193][0] ),
    .C(_09539_),
    .X(_10068_));
 sky130_fd_sc_hd__nand2_8 _14343_ (.A(_09673_),
    .B(_08994_),
    .Y(_10069_));
 sky130_fd_sc_hd__inv_2 _14344_ (.A(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__buf_4 _14345_ (.A(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__and3_1 _14346_ (.A(_10071_),
    .B(\line_cache[192][0] ),
    .C(_09539_),
    .X(_10072_));
 sky130_fd_sc_hd__nand2_8 _14347_ (.A(_09558_),
    .B(_09778_),
    .Y(_10073_));
 sky130_fd_sc_hd__inv_4 _14348_ (.A(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__clkbuf_4 _14349_ (.A(_09538_),
    .X(_10075_));
 sky130_fd_sc_hd__and3_1 _14350_ (.A(_10074_),
    .B(\line_cache[194][0] ),
    .C(_10075_),
    .X(_10076_));
 sky130_fd_sc_hd__a2111o_1 _14351_ (.A1(_10066_),
    .A2(\line_cache[286][0] ),
    .B1(_10068_),
    .C1(_10072_),
    .D1(_10076_),
    .X(_10077_));
 sky130_fd_sc_hd__or4_1 _14352_ (.A(_10043_),
    .B(_10053_),
    .C(_10065_),
    .D(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__a22o_1 _14353_ (.A1(_09623_),
    .A2(\line_cache[275][0] ),
    .B1(_09620_),
    .B2(\line_cache[274][0] ),
    .X(_10079_));
 sky130_fd_sc_hd__inv_2 _14354_ (.A(_09630_),
    .Y(_10080_));
 sky130_fd_sc_hd__inv_2 _14355_ (.A(_09632_),
    .Y(_10081_));
 sky130_fd_sc_hd__a22o_1 _14356_ (.A1(_10080_),
    .A2(\line_cache[276][0] ),
    .B1(\line_cache[277][0] ),
    .B2(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__inv_2 _14357_ (.A(_09625_),
    .Y(_10083_));
 sky130_fd_sc_hd__inv_2 _14358_ (.A(_09627_),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(_09868_),
    .B(_09551_),
    .Y(_10085_));
 sky130_fd_sc_hd__inv_2 _14360_ (.A(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_1 _14361_ (.A(_09871_),
    .B(_09551_),
    .Y(_10087_));
 sky130_fd_sc_hd__inv_2 _14362_ (.A(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__a22o_1 _14363_ (.A1(_10086_),
    .A2(\line_cache[270][0] ),
    .B1(\line_cache[269][0] ),
    .B2(_10088_),
    .X(_10089_));
 sky130_fd_sc_hd__a221o_1 _14364_ (.A1(\line_cache[273][0] ),
    .A2(_10083_),
    .B1(\line_cache[272][0] ),
    .B2(_10084_),
    .C1(_10089_),
    .X(_10090_));
 sky130_fd_sc_hd__a22o_1 _14365_ (.A1(_09663_),
    .A2(\line_cache[281][0] ),
    .B1(\line_cache[280][0] ),
    .B2(_09655_),
    .X(_10091_));
 sky130_fd_sc_hd__a22oi_1 _14366_ (.A1(_09661_),
    .A2(\line_cache[282][0] ),
    .B1(\line_cache[283][0] ),
    .B2(_09658_),
    .Y(_10092_));
 sky130_fd_sc_hd__a22oi_1 _14367_ (.A1(_09645_),
    .A2(\line_cache[285][0] ),
    .B1(\line_cache[284][0] ),
    .B2(_09648_),
    .Y(_10093_));
 sky130_fd_sc_hd__a22oi_1 _14368_ (.A1(_09636_),
    .A2(\line_cache[278][0] ),
    .B1(\line_cache[279][0] ),
    .B2(_09639_),
    .Y(_10094_));
 sky130_fd_sc_hd__and4b_1 _14369_ (.A_N(_10091_),
    .B(_10092_),
    .C(_10093_),
    .D(_10094_),
    .X(_10095_));
 sky130_fd_sc_hd__or4b_2 _14370_ (.A(_10079_),
    .B(_10082_),
    .C(_10090_),
    .D_N(_10095_),
    .X(_10096_));
 sky130_fd_sc_hd__nor2_1 _14371_ (.A(_10078_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__buf_6 _14372_ (.A(_09595_),
    .X(_10098_));
 sky130_fd_sc_hd__clkinv_4 _14373_ (.A(_09550_),
    .Y(_10099_));
 sky130_fd_sc_hd__clkbuf_4 _14374_ (.A(_10099_),
    .X(_10100_));
 sky130_fd_sc_hd__and3_1 _14375_ (.A(_10098_),
    .B(\line_cache[229][0] ),
    .C(_10100_),
    .X(_10101_));
 sky130_fd_sc_hd__buf_8 _14376_ (.A(_10044_),
    .X(_10102_));
 sky130_fd_sc_hd__and3_1 _14377_ (.A(_10102_),
    .B(\line_cache[230][0] ),
    .C(_10100_),
    .X(_10103_));
 sky130_fd_sc_hd__clkinv_4 _14378_ (.A(_10048_),
    .Y(_10104_));
 sky130_fd_sc_hd__and3_1 _14379_ (.A(_10104_),
    .B(\line_cache[227][0] ),
    .C(_10100_),
    .X(_10105_));
 sky130_fd_sc_hd__inv_4 _14380_ (.A(_10050_),
    .Y(_10106_));
 sky130_fd_sc_hd__and3_1 _14381_ (.A(_10106_),
    .B(\line_cache[228][0] ),
    .C(_10100_),
    .X(_10107_));
 sky130_fd_sc_hd__or4_1 _14382_ (.A(_10101_),
    .B(_10103_),
    .C(_10105_),
    .D(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__buf_8 _14383_ (.A(_09600_),
    .X(_10109_));
 sky130_fd_sc_hd__and3_1 _14384_ (.A(_09544_),
    .B(\line_cache[223][0] ),
    .C(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__and3_1 _14385_ (.A(_10071_),
    .B(\line_cache[224][0] ),
    .C(_10100_),
    .X(_10111_));
 sky130_fd_sc_hd__and3_1 _14386_ (.A(_10067_),
    .B(\line_cache[225][0] ),
    .C(_10100_),
    .X(_10112_));
 sky130_fd_sc_hd__and3_1 _14387_ (.A(_10074_),
    .B(\line_cache[226][0] ),
    .C(_10100_),
    .X(_10113_));
 sky130_fd_sc_hd__or4_1 _14388_ (.A(_10110_),
    .B(_10111_),
    .C(_10112_),
    .D(_10113_),
    .X(_10114_));
 sky130_fd_sc_hd__inv_12 _14389_ (.A(_10037_),
    .Y(_10115_));
 sky130_fd_sc_hd__nor2_2 _14390_ (.A(_09550_),
    .B(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__nor2_2 _14391_ (.A(_09550_),
    .B(_10032_),
    .Y(_10117_));
 sky130_fd_sc_hd__nor2_2 _14392_ (.A(_09550_),
    .B(_10040_),
    .Y(_10118_));
 sky130_fd_sc_hd__clkinv_16 _14393_ (.A(_10034_),
    .Y(_10119_));
 sky130_fd_sc_hd__nor2_2 _14394_ (.A(_09550_),
    .B(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__a22o_1 _14395_ (.A1(_10118_),
    .A2(\line_cache[236][0] ),
    .B1(_10120_),
    .B2(\line_cache[235][0] ),
    .X(_10121_));
 sky130_fd_sc_hd__a221o_1 _14396_ (.A1(\line_cache[238][0] ),
    .A2(_10116_),
    .B1(\line_cache[237][0] ),
    .B2(_10117_),
    .C1(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__nor2_2 _14397_ (.A(_09550_),
    .B(_10055_),
    .Y(_10123_));
 sky130_fd_sc_hd__nor2_2 _14398_ (.A(_09550_),
    .B(_10058_),
    .Y(_10124_));
 sky130_fd_sc_hd__nor2_4 _14399_ (.A(_09550_),
    .B(_09578_),
    .Y(_10125_));
 sky130_fd_sc_hd__nor2_4 _14400_ (.A(_09550_),
    .B(_10062_),
    .Y(_10126_));
 sky130_fd_sc_hd__a22o_1 _14401_ (.A1(_10125_),
    .A2(\line_cache[232][0] ),
    .B1(_10126_),
    .B2(\line_cache[231][0] ),
    .X(_10127_));
 sky130_fd_sc_hd__a221o_1 _14402_ (.A1(\line_cache[234][0] ),
    .A2(_10123_),
    .B1(\line_cache[233][0] ),
    .B2(_10124_),
    .C1(_10127_),
    .X(_10128_));
 sky130_fd_sc_hd__or4_1 _14403_ (.A(_10108_),
    .B(_10114_),
    .C(_10122_),
    .D(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__nor2_2 _14404_ (.A(_09543_),
    .B(_10115_),
    .Y(_10130_));
 sky130_fd_sc_hd__nor2_2 _14405_ (.A(_09543_),
    .B(_10032_),
    .Y(_10131_));
 sky130_fd_sc_hd__nor2_2 _14406_ (.A(_09543_),
    .B(_10040_),
    .Y(_10132_));
 sky130_fd_sc_hd__nor2_2 _14407_ (.A(_09543_),
    .B(_10119_),
    .Y(_10133_));
 sky130_fd_sc_hd__a22o_1 _14408_ (.A1(_10132_),
    .A2(\line_cache[220][0] ),
    .B1(_10133_),
    .B2(\line_cache[219][0] ),
    .X(_10134_));
 sky130_fd_sc_hd__a221o_1 _14409_ (.A1(\line_cache[222][0] ),
    .A2(_10130_),
    .B1(\line_cache[221][0] ),
    .B2(_10131_),
    .C1(_10134_),
    .X(_10135_));
 sky130_fd_sc_hd__nor2_2 _14410_ (.A(_09543_),
    .B(_10073_),
    .Y(_10136_));
 sky130_fd_sc_hd__nor2_4 _14411_ (.A(_09543_),
    .B(_09569_),
    .Y(_10137_));
 sky130_fd_sc_hd__nor2_4 _14412_ (.A(_09543_),
    .B(_10069_),
    .Y(_10138_));
 sky130_fd_sc_hd__and3_4 _14413_ (.A(_09538_),
    .B(_09616_),
    .C(_10109_),
    .X(_10139_));
 sky130_fd_sc_hd__a22o_1 _14414_ (.A1(_10138_),
    .A2(\line_cache[208][0] ),
    .B1(_10139_),
    .B2(\line_cache[207][0] ),
    .X(_10140_));
 sky130_fd_sc_hd__a221o_1 _14415_ (.A1(\line_cache[210][0] ),
    .A2(_10136_),
    .B1(\line_cache[209][0] ),
    .B2(_10137_),
    .C1(_10140_),
    .X(_10141_));
 sky130_fd_sc_hd__nor2_2 _14416_ (.A(_09543_),
    .B(_10055_),
    .Y(_10142_));
 sky130_fd_sc_hd__nor2_2 _14417_ (.A(_09543_),
    .B(_10058_),
    .Y(_10143_));
 sky130_fd_sc_hd__nor2_2 _14418_ (.A(_09543_),
    .B(_09578_),
    .Y(_10144_));
 sky130_fd_sc_hd__nor2_2 _14419_ (.A(_09543_),
    .B(_10062_),
    .Y(_10145_));
 sky130_fd_sc_hd__a22o_1 _14420_ (.A1(_10144_),
    .A2(\line_cache[216][0] ),
    .B1(_10145_),
    .B2(\line_cache[215][0] ),
    .X(_10146_));
 sky130_fd_sc_hd__a221o_1 _14421_ (.A1(\line_cache[218][0] ),
    .A2(_10142_),
    .B1(\line_cache[217][0] ),
    .B2(_10143_),
    .C1(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__or2_2 _14422_ (.A(_09543_),
    .B(_10048_),
    .X(_10148_));
 sky130_fd_sc_hd__and2b_1 _14423_ (.A_N(_10148_),
    .B(\line_cache[211][0] ),
    .X(_10149_));
 sky130_fd_sc_hd__or2_2 _14424_ (.A(_09543_),
    .B(_10050_),
    .X(_10150_));
 sky130_fd_sc_hd__and2b_1 _14425_ (.A_N(_10150_),
    .B(\line_cache[212][0] ),
    .X(_10151_));
 sky130_fd_sc_hd__or2_2 _14426_ (.A(_09543_),
    .B(_09596_),
    .X(_10152_));
 sky130_fd_sc_hd__and2b_1 _14427_ (.A_N(_10152_),
    .B(\line_cache[213][0] ),
    .X(_10153_));
 sky130_fd_sc_hd__or2_2 _14428_ (.A(_09543_),
    .B(_10045_),
    .X(_10154_));
 sky130_fd_sc_hd__and2b_1 _14429_ (.A_N(_10154_),
    .B(\line_cache[214][0] ),
    .X(_10155_));
 sky130_fd_sc_hd__or4_1 _14430_ (.A(_10149_),
    .B(_10151_),
    .C(_10153_),
    .D(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__or4_2 _14431_ (.A(_10135_),
    .B(_10141_),
    .C(_10147_),
    .D(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__nor2_1 _14432_ (.A(_10129_),
    .B(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__nor2_4 _14433_ (.A(_09766_),
    .B(_10062_),
    .Y(_10159_));
 sky130_fd_sc_hd__inv_2 _14434_ (.A(_09766_),
    .Y(_10160_));
 sky130_fd_sc_hd__buf_4 _14435_ (.A(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__and3_1 _14436_ (.A(_10102_),
    .B(\line_cache[70][0] ),
    .C(_10161_),
    .X(_10162_));
 sky130_fd_sc_hd__nor2_4 _14437_ (.A(_09766_),
    .B(_10050_),
    .Y(_10163_));
 sky130_fd_sc_hd__nor2_4 _14438_ (.A(_09766_),
    .B(_09596_),
    .Y(_10164_));
 sky130_fd_sc_hd__a22o_1 _14439_ (.A1(_10163_),
    .A2(\line_cache[68][0] ),
    .B1(_10164_),
    .B2(\line_cache[69][0] ),
    .X(_10165_));
 sky130_fd_sc_hd__a211o_1 _14440_ (.A1(\line_cache[71][0] ),
    .A2(_10159_),
    .B1(_10162_),
    .C1(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__buf_4 _14441_ (.A(_10160_),
    .X(_10167_));
 sky130_fd_sc_hd__and3_2 _14442_ (.A(_10167_),
    .B(_09531_),
    .C(_10109_),
    .X(_10168_));
 sky130_fd_sc_hd__and3_1 _14443_ (.A(_10031_),
    .B(\line_cache[77][0] ),
    .C(_10161_),
    .X(_10169_));
 sky130_fd_sc_hd__and3_1 _14444_ (.A(_10038_),
    .B(\line_cache[78][0] ),
    .C(_10161_),
    .X(_10170_));
 sky130_fd_sc_hd__and3_1 _14445_ (.A(_10041_),
    .B(\line_cache[76][0] ),
    .C(_10161_),
    .X(_10171_));
 sky130_fd_sc_hd__a2111o_1 _14446_ (.A1(_10168_),
    .A2(\line_cache[79][0] ),
    .B1(_10169_),
    .C1(_10170_),
    .D1(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__nor2_4 _14447_ (.A(_09766_),
    .B(_10119_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor2_4 _14448_ (.A(_09766_),
    .B(_10055_),
    .Y(_10174_));
 sky130_fd_sc_hd__nor2_4 _14449_ (.A(_09766_),
    .B(_09578_),
    .Y(_10175_));
 sky130_fd_sc_hd__clkbuf_8 _14450_ (.A(_10057_),
    .X(_10176_));
 sky130_fd_sc_hd__and3_1 _14451_ (.A(_10176_),
    .B(\line_cache[73][0] ),
    .C(_10161_),
    .X(_10177_));
 sky130_fd_sc_hd__a21o_1 _14452_ (.A1(\line_cache[72][0] ),
    .A2(_10175_),
    .B1(_10177_),
    .X(_10178_));
 sky130_fd_sc_hd__a221o_1 _14453_ (.A1(\line_cache[75][0] ),
    .A2(_10173_),
    .B1(\line_cache[74][0] ),
    .B2(_10174_),
    .C1(_10178_),
    .X(_10179_));
 sky130_fd_sc_hd__nor2_4 _14454_ (.A(_09766_),
    .B(_10048_),
    .Y(_10180_));
 sky130_fd_sc_hd__nor2_4 _14455_ (.A(_09766_),
    .B(_10073_),
    .Y(_10181_));
 sky130_fd_sc_hd__nor2_4 _14456_ (.A(_09766_),
    .B(_10069_),
    .Y(_10182_));
 sky130_fd_sc_hd__nor2_4 _14457_ (.A(_09766_),
    .B(_09569_),
    .Y(_10183_));
 sky130_fd_sc_hd__a22o_1 _14458_ (.A1(_10182_),
    .A2(\line_cache[64][0] ),
    .B1(_10183_),
    .B2(\line_cache[65][0] ),
    .X(_10184_));
 sky130_fd_sc_hd__a221o_1 _14459_ (.A1(\line_cache[67][0] ),
    .A2(_10180_),
    .B1(\line_cache[66][0] ),
    .B2(_10181_),
    .C1(_10184_),
    .X(_10185_));
 sky130_fd_sc_hd__or4_4 _14460_ (.A(_10166_),
    .B(_10172_),
    .C(_10179_),
    .D(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__nor2_2 _14461_ (.A(_09555_),
    .B(_10115_),
    .Y(_10187_));
 sky130_fd_sc_hd__nor2_2 _14462_ (.A(_09555_),
    .B(_10032_),
    .Y(_10188_));
 sky130_fd_sc_hd__nor2_2 _14463_ (.A(_09555_),
    .B(_10040_),
    .Y(_10189_));
 sky130_fd_sc_hd__nor2_2 _14464_ (.A(_09555_),
    .B(_10119_),
    .Y(_10190_));
 sky130_fd_sc_hd__a22o_1 _14465_ (.A1(_10189_),
    .A2(\line_cache[252][0] ),
    .B1(_10190_),
    .B2(\line_cache[251][0] ),
    .X(_10191_));
 sky130_fd_sc_hd__a221o_1 _14466_ (.A1(\line_cache[254][0] ),
    .A2(_10187_),
    .B1(\line_cache[253][0] ),
    .B2(_10188_),
    .C1(_10191_),
    .X(_10192_));
 sky130_fd_sc_hd__nor2_2 _14467_ (.A(_09555_),
    .B(_10055_),
    .Y(_10193_));
 sky130_fd_sc_hd__nor2_2 _14468_ (.A(_09555_),
    .B(_10058_),
    .Y(_10194_));
 sky130_fd_sc_hd__nor2_2 _14469_ (.A(_09555_),
    .B(_09578_),
    .Y(_10195_));
 sky130_fd_sc_hd__nor2_2 _14470_ (.A(_09555_),
    .B(_10062_),
    .Y(_10196_));
 sky130_fd_sc_hd__a22o_1 _14471_ (.A1(_10195_),
    .A2(\line_cache[248][0] ),
    .B1(_10196_),
    .B2(\line_cache[247][0] ),
    .X(_10197_));
 sky130_fd_sc_hd__a221o_1 _14472_ (.A1(\line_cache[250][0] ),
    .A2(_10193_),
    .B1(\line_cache[249][0] ),
    .B2(_10194_),
    .C1(_10197_),
    .X(_10198_));
 sky130_fd_sc_hd__and3_2 _14473_ (.A(_10100_),
    .B(_09531_),
    .C(_10109_),
    .X(_10199_));
 sky130_fd_sc_hd__or2_2 _14474_ (.A(_09554_),
    .B(_10069_),
    .X(_10200_));
 sky130_fd_sc_hd__and2b_1 _14475_ (.A_N(_10200_),
    .B(\line_cache[240][0] ),
    .X(_10201_));
 sky130_fd_sc_hd__and2b_1 _14476_ (.A_N(_09570_),
    .B(\line_cache[241][0] ),
    .X(_10202_));
 sky130_fd_sc_hd__or2_2 _14477_ (.A(_09554_),
    .B(_10073_),
    .X(_10203_));
 sky130_fd_sc_hd__and2b_1 _14478_ (.A_N(_10203_),
    .B(\line_cache[242][0] ),
    .X(_10204_));
 sky130_fd_sc_hd__a2111o_1 _14479_ (.A1(\line_cache[239][0] ),
    .A2(_10199_),
    .B1(_10201_),
    .C1(_10202_),
    .D1(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__or2_2 _14480_ (.A(_09554_),
    .B(_10048_),
    .X(_10206_));
 sky130_fd_sc_hd__and2b_1 _14481_ (.A_N(_10206_),
    .B(\line_cache[243][0] ),
    .X(_10207_));
 sky130_fd_sc_hd__or2_2 _14482_ (.A(_09554_),
    .B(_10050_),
    .X(_10208_));
 sky130_fd_sc_hd__and2b_1 _14483_ (.A_N(_10208_),
    .B(\line_cache[244][0] ),
    .X(_10209_));
 sky130_fd_sc_hd__and2b_1 _14484_ (.A_N(_09597_),
    .B(\line_cache[245][0] ),
    .X(_10210_));
 sky130_fd_sc_hd__or2_2 _14485_ (.A(_09554_),
    .B(_10045_),
    .X(_10211_));
 sky130_fd_sc_hd__and2b_1 _14486_ (.A_N(_10211_),
    .B(\line_cache[246][0] ),
    .X(_10212_));
 sky130_fd_sc_hd__or4_1 _14487_ (.A(_10207_),
    .B(_10209_),
    .C(_10210_),
    .D(_10212_),
    .X(_10213_));
 sky130_fd_sc_hd__or4_1 _14488_ (.A(_10192_),
    .B(_10198_),
    .C(_10205_),
    .D(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__nor2_1 _14489_ (.A(_10186_),
    .B(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__and4_2 _14490_ (.A(_10030_),
    .B(_10097_),
    .C(_10158_),
    .D(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__and3_4 _14491_ (.A(_09753_),
    .B(_09531_),
    .C(_10109_),
    .X(_10217_));
 sky130_fd_sc_hd__nor2_4 _14492_ (.A(_10115_),
    .B(_09754_),
    .Y(_10218_));
 sky130_fd_sc_hd__nor2_4 _14493_ (.A(_10032_),
    .B(_09754_),
    .Y(_10219_));
 sky130_fd_sc_hd__nor2_4 _14494_ (.A(_10040_),
    .B(_09754_),
    .Y(_10220_));
 sky130_fd_sc_hd__a22o_1 _14495_ (.A1(_10219_),
    .A2(\line_cache[157][0] ),
    .B1(\line_cache[156][0] ),
    .B2(_10220_),
    .X(_10221_));
 sky130_fd_sc_hd__a221o_1 _14496_ (.A1(\line_cache[159][0] ),
    .A2(_10217_),
    .B1(\line_cache[158][0] ),
    .B2(_10218_),
    .C1(_10221_),
    .X(_10222_));
 sky130_fd_sc_hd__nor2_4 _14497_ (.A(_09596_),
    .B(_09754_),
    .Y(_10223_));
 sky130_fd_sc_hd__nor2_4 _14498_ (.A(_10050_),
    .B(_09754_),
    .Y(_10224_));
 sky130_fd_sc_hd__nor2_4 _14499_ (.A(_10062_),
    .B(_09754_),
    .Y(_10225_));
 sky130_fd_sc_hd__nor2_4 _14500_ (.A(_10045_),
    .B(_09754_),
    .Y(_10226_));
 sky130_fd_sc_hd__a22o_1 _14501_ (.A1(_10225_),
    .A2(\line_cache[151][0] ),
    .B1(\line_cache[150][0] ),
    .B2(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__a221oi_2 _14502_ (.A1(\line_cache[149][0] ),
    .A2(_10223_),
    .B1(\line_cache[148][0] ),
    .B2(_10224_),
    .C1(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__nor2_4 _14503_ (.A(_09569_),
    .B(_09754_),
    .Y(_10229_));
 sky130_fd_sc_hd__nor2_4 _14504_ (.A(_10069_),
    .B(_09754_),
    .Y(_10230_));
 sky130_fd_sc_hd__nor2_4 _14505_ (.A(_10048_),
    .B(_09754_),
    .Y(_10231_));
 sky130_fd_sc_hd__nor2_4 _14506_ (.A(_10073_),
    .B(_09754_),
    .Y(_10232_));
 sky130_fd_sc_hd__a22o_1 _14507_ (.A1(_10231_),
    .A2(\line_cache[147][0] ),
    .B1(\line_cache[146][0] ),
    .B2(_10232_),
    .X(_10233_));
 sky130_fd_sc_hd__a221oi_1 _14508_ (.A1(\line_cache[145][0] ),
    .A2(_10229_),
    .B1(\line_cache[144][0] ),
    .B2(_10230_),
    .C1(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__nor2_4 _14509_ (.A(_10058_),
    .B(_09754_),
    .Y(_10235_));
 sky130_fd_sc_hd__nor2_4 _14510_ (.A(_09578_),
    .B(_09754_),
    .Y(_10236_));
 sky130_fd_sc_hd__nor2_4 _14511_ (.A(_10119_),
    .B(_09754_),
    .Y(_10237_));
 sky130_fd_sc_hd__nor2_4 _14512_ (.A(_10055_),
    .B(_09754_),
    .Y(_10238_));
 sky130_fd_sc_hd__a22o_1 _14513_ (.A1(_10237_),
    .A2(\line_cache[155][0] ),
    .B1(\line_cache[154][0] ),
    .B2(_10238_),
    .X(_10239_));
 sky130_fd_sc_hd__a221oi_2 _14514_ (.A1(\line_cache[153][0] ),
    .A2(_10235_),
    .B1(\line_cache[152][0] ),
    .B2(_10236_),
    .C1(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__and4b_1 _14515_ (.A_N(_10222_),
    .B(_10228_),
    .C(_10234_),
    .D(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__and3_4 _14516_ (.A(_09751_),
    .B(_09531_),
    .C(_10109_),
    .X(_10242_));
 sky130_fd_sc_hd__nor2_4 _14517_ (.A(_10115_),
    .B(_09752_),
    .Y(_10243_));
 sky130_fd_sc_hd__nor2_4 _14518_ (.A(_10032_),
    .B(_09752_),
    .Y(_10244_));
 sky130_fd_sc_hd__nor2_4 _14519_ (.A(_10040_),
    .B(_09752_),
    .Y(_10245_));
 sky130_fd_sc_hd__a22o_1 _14520_ (.A1(_10244_),
    .A2(\line_cache[173][0] ),
    .B1(\line_cache[172][0] ),
    .B2(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__a221o_1 _14521_ (.A1(\line_cache[175][0] ),
    .A2(_10242_),
    .B1(\line_cache[174][0] ),
    .B2(_10243_),
    .C1(_10246_),
    .X(_10247_));
 sky130_fd_sc_hd__nor2_2 _14522_ (.A(_10062_),
    .B(_09752_),
    .Y(_10248_));
 sky130_fd_sc_hd__nor2_2 _14523_ (.A(_10045_),
    .B(_09752_),
    .Y(_10249_));
 sky130_fd_sc_hd__nor2_2 _14524_ (.A(_09596_),
    .B(_09752_),
    .Y(_10250_));
 sky130_fd_sc_hd__nor2_2 _14525_ (.A(_10050_),
    .B(_09752_),
    .Y(_10251_));
 sky130_fd_sc_hd__a22o_1 _14526_ (.A1(_10250_),
    .A2(\line_cache[165][0] ),
    .B1(\line_cache[164][0] ),
    .B2(_10251_),
    .X(_10252_));
 sky130_fd_sc_hd__a221oi_1 _14527_ (.A1(\line_cache[167][0] ),
    .A2(_10248_),
    .B1(\line_cache[166][0] ),
    .B2(_10249_),
    .C1(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__nor2_2 _14528_ (.A(_10048_),
    .B(_09752_),
    .Y(_10254_));
 sky130_fd_sc_hd__nor2_4 _14529_ (.A(_10073_),
    .B(_09752_),
    .Y(_10255_));
 sky130_fd_sc_hd__nor2_4 _14530_ (.A(_10069_),
    .B(_09752_),
    .Y(_10256_));
 sky130_fd_sc_hd__nor2_4 _14531_ (.A(_09569_),
    .B(_09752_),
    .Y(_10257_));
 sky130_fd_sc_hd__a22o_1 _14532_ (.A1(_10256_),
    .A2(\line_cache[160][0] ),
    .B1(\line_cache[161][0] ),
    .B2(_10257_),
    .X(_10258_));
 sky130_fd_sc_hd__a221oi_2 _14533_ (.A1(\line_cache[163][0] ),
    .A2(_10254_),
    .B1(\line_cache[162][0] ),
    .B2(_10255_),
    .C1(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__nor2_4 _14534_ (.A(_10058_),
    .B(_09752_),
    .Y(_10260_));
 sky130_fd_sc_hd__nor2_4 _14535_ (.A(_09578_),
    .B(_09752_),
    .Y(_10261_));
 sky130_fd_sc_hd__nor2_4 _14536_ (.A(_10119_),
    .B(_09752_),
    .Y(_10262_));
 sky130_fd_sc_hd__nor2_4 _14537_ (.A(_10055_),
    .B(_09752_),
    .Y(_10263_));
 sky130_fd_sc_hd__a22o_1 _14538_ (.A1(_10262_),
    .A2(\line_cache[171][0] ),
    .B1(\line_cache[170][0] ),
    .B2(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__a221oi_2 _14539_ (.A1(\line_cache[169][0] ),
    .A2(_10260_),
    .B1(\line_cache[168][0] ),
    .B2(_10261_),
    .C1(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__and4b_1 _14540_ (.A_N(_10247_),
    .B(_10253_),
    .C(_10259_),
    .D(_10265_),
    .X(_10266_));
 sky130_fd_sc_hd__nor2_2 _14541_ (.A(_09551_),
    .B(_09601_),
    .Y(_10267_));
 sky130_fd_sc_hd__inv_2 _14542_ (.A(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__nor2_4 _14543_ (.A(_10268_),
    .B(_09756_),
    .Y(_10269_));
 sky130_fd_sc_hd__nor2_4 _14544_ (.A(_09756_),
    .B(_10115_),
    .Y(_10270_));
 sky130_fd_sc_hd__nor2_4 _14545_ (.A(_10040_),
    .B(_09756_),
    .Y(_10271_));
 sky130_fd_sc_hd__nor2_4 _14546_ (.A(_10032_),
    .B(_09756_),
    .Y(_10272_));
 sky130_fd_sc_hd__a22o_1 _14547_ (.A1(_10271_),
    .A2(\line_cache[188][0] ),
    .B1(\line_cache[189][0] ),
    .B2(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__a221oi_1 _14548_ (.A1(\line_cache[191][0] ),
    .A2(_10269_),
    .B1(\line_cache[190][0] ),
    .B2(_10270_),
    .C1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__nor2_4 _14549_ (.A(_10119_),
    .B(_09756_),
    .Y(_10275_));
 sky130_fd_sc_hd__nor2_4 _14550_ (.A(_09756_),
    .B(_10055_),
    .Y(_10276_));
 sky130_fd_sc_hd__nor2_4 _14551_ (.A(_09578_),
    .B(_09756_),
    .Y(_10277_));
 sky130_fd_sc_hd__nor2_4 _14552_ (.A(_10058_),
    .B(_09756_),
    .Y(_10278_));
 sky130_fd_sc_hd__a22o_1 _14553_ (.A1(_10277_),
    .A2(\line_cache[184][0] ),
    .B1(\line_cache[185][0] ),
    .B2(_10278_),
    .X(_10279_));
 sky130_fd_sc_hd__a221oi_4 _14554_ (.A1(\line_cache[187][0] ),
    .A2(_10275_),
    .B1(\line_cache[186][0] ),
    .B2(_10276_),
    .C1(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__nand2_1 _14555_ (.A(_10274_),
    .B(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__nor2_4 _14556_ (.A(_10048_),
    .B(_09756_),
    .Y(_10282_));
 sky130_fd_sc_hd__nor2_4 _14557_ (.A(_10073_),
    .B(_09756_),
    .Y(_10283_));
 sky130_fd_sc_hd__nor2_2 _14558_ (.A(_10069_),
    .B(_09756_),
    .Y(_10284_));
 sky130_fd_sc_hd__nor2_4 _14559_ (.A(_09569_),
    .B(_09756_),
    .Y(_10285_));
 sky130_fd_sc_hd__a22o_1 _14560_ (.A1(_10284_),
    .A2(\line_cache[176][0] ),
    .B1(_10285_),
    .B2(\line_cache[177][0] ),
    .X(_10286_));
 sky130_fd_sc_hd__a221o_1 _14561_ (.A1(\line_cache[179][0] ),
    .A2(_10282_),
    .B1(\line_cache[178][0] ),
    .B2(_10283_),
    .C1(_10286_),
    .X(_10287_));
 sky130_fd_sc_hd__buf_4 _14562_ (.A(_09755_),
    .X(_10288_));
 sky130_fd_sc_hd__clkbuf_8 _14563_ (.A(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__and3_1 _14564_ (.A(_10289_),
    .B(_10098_),
    .C(\line_cache[181][0] ),
    .X(_10290_));
 sky130_fd_sc_hd__and3_1 _14565_ (.A(_10288_),
    .B(\line_cache[183][0] ),
    .C(_10061_),
    .X(_10291_));
 sky130_fd_sc_hd__a31o_1 _14566_ (.A1(\line_cache[182][0] ),
    .A2(_10289_),
    .A3(_10102_),
    .B1(_10291_),
    .X(_10292_));
 sky130_fd_sc_hd__a311o_1 _14567_ (.A1(\line_cache[180][0] ),
    .A2(_10289_),
    .A3(_10106_),
    .B1(_10290_),
    .C1(_10292_),
    .X(_10293_));
 sky130_fd_sc_hd__nor3_1 _14568_ (.A(_10281_),
    .B(_10287_),
    .C(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__and3_2 _14569_ (.A(_10241_),
    .B(_10266_),
    .C(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__nor2_4 _14570_ (.A(_09768_),
    .B(_10048_),
    .Y(_10296_));
 sky130_fd_sc_hd__nor2_4 _14571_ (.A(_09768_),
    .B(_10073_),
    .Y(_10297_));
 sky130_fd_sc_hd__nor2_2 _14572_ (.A(_09768_),
    .B(_10069_),
    .Y(_10298_));
 sky130_fd_sc_hd__nor2_2 _14573_ (.A(_09768_),
    .B(_09569_),
    .Y(_10299_));
 sky130_fd_sc_hd__a22o_1 _14574_ (.A1(_10298_),
    .A2(\line_cache[112][0] ),
    .B1(_10299_),
    .B2(\line_cache[113][0] ),
    .X(_10300_));
 sky130_fd_sc_hd__a221o_1 _14575_ (.A1(\line_cache[115][0] ),
    .A2(_10296_),
    .B1(\line_cache[114][0] ),
    .B2(_10297_),
    .C1(_10300_),
    .X(_10301_));
 sky130_fd_sc_hd__inv_2 _14576_ (.A(_09767_),
    .Y(_10302_));
 sky130_fd_sc_hd__and3_1 _14577_ (.A(_10302_),
    .B(_09531_),
    .C(_10109_),
    .X(_10303_));
 sky130_fd_sc_hd__nor2_2 _14578_ (.A(_09768_),
    .B(_10115_),
    .Y(_10304_));
 sky130_fd_sc_hd__nor2_2 _14579_ (.A(_09768_),
    .B(_10040_),
    .Y(_10305_));
 sky130_fd_sc_hd__nor2_2 _14580_ (.A(_09768_),
    .B(_10032_),
    .Y(_10306_));
 sky130_fd_sc_hd__a22o_1 _14581_ (.A1(_10305_),
    .A2(\line_cache[124][0] ),
    .B1(_10306_),
    .B2(\line_cache[125][0] ),
    .X(_10307_));
 sky130_fd_sc_hd__a221o_1 _14582_ (.A1(\line_cache[127][0] ),
    .A2(_10303_),
    .B1(\line_cache[126][0] ),
    .B2(_10304_),
    .C1(_10307_),
    .X(_10308_));
 sky130_fd_sc_hd__nor2_2 _14583_ (.A(_09768_),
    .B(_10062_),
    .Y(_10309_));
 sky130_fd_sc_hd__nor2_2 _14584_ (.A(_09768_),
    .B(_10045_),
    .Y(_10310_));
 sky130_fd_sc_hd__nor2_4 _14585_ (.A(_09768_),
    .B(_10050_),
    .Y(_10311_));
 sky130_fd_sc_hd__nor2_4 _14586_ (.A(_09768_),
    .B(_09596_),
    .Y(_10312_));
 sky130_fd_sc_hd__a22o_1 _14587_ (.A1(_10311_),
    .A2(\line_cache[116][0] ),
    .B1(_10312_),
    .B2(\line_cache[117][0] ),
    .X(_10313_));
 sky130_fd_sc_hd__a221o_1 _14588_ (.A1(\line_cache[119][0] ),
    .A2(_10309_),
    .B1(\line_cache[118][0] ),
    .B2(_10310_),
    .C1(_10313_),
    .X(_10314_));
 sky130_fd_sc_hd__nor2_4 _14589_ (.A(_09768_),
    .B(_10119_),
    .Y(_10315_));
 sky130_fd_sc_hd__nor2_4 _14590_ (.A(_09768_),
    .B(_10055_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_4 _14591_ (.A(_09768_),
    .B(_09578_),
    .Y(_10317_));
 sky130_fd_sc_hd__nor2_1 _14592_ (.A(_09768_),
    .B(_10058_),
    .Y(_10318_));
 sky130_fd_sc_hd__a22o_1 _14593_ (.A1(_10317_),
    .A2(\line_cache[120][0] ),
    .B1(_10318_),
    .B2(\line_cache[121][0] ),
    .X(_10319_));
 sky130_fd_sc_hd__a221o_1 _14594_ (.A1(\line_cache[123][0] ),
    .A2(_10315_),
    .B1(\line_cache[122][0] ),
    .B2(_10316_),
    .C1(_10319_),
    .X(_10320_));
 sky130_fd_sc_hd__or4_1 _14595_ (.A(_10301_),
    .B(_10308_),
    .C(_10314_),
    .D(_10320_),
    .X(_10321_));
 sky130_fd_sc_hd__nor2_4 _14596_ (.A(_10062_),
    .B(_09760_),
    .Y(_10322_));
 sky130_fd_sc_hd__nor2_4 _14597_ (.A(_09760_),
    .B(_10045_),
    .Y(_10323_));
 sky130_fd_sc_hd__nor2_4 _14598_ (.A(_10050_),
    .B(_09759_),
    .Y(_10324_));
 sky130_fd_sc_hd__and3_1 _14599_ (.A(_09758_),
    .B(_10098_),
    .C(\line_cache[133][0] ),
    .X(_10325_));
 sky130_fd_sc_hd__a21o_1 _14600_ (.A1(\line_cache[132][0] ),
    .A2(_10324_),
    .B1(_10325_),
    .X(_10326_));
 sky130_fd_sc_hd__a221o_1 _14601_ (.A1(\line_cache[135][0] ),
    .A2(_10322_),
    .B1(\line_cache[134][0] ),
    .B2(_10323_),
    .C1(_10326_),
    .X(_10327_));
 sky130_fd_sc_hd__nor2_2 _14602_ (.A(_10048_),
    .B(_09760_),
    .Y(_10328_));
 sky130_fd_sc_hd__nor2_2 _14603_ (.A(_09760_),
    .B(_10073_),
    .Y(_10329_));
 sky130_fd_sc_hd__nor2_2 _14604_ (.A(_09569_),
    .B(_09760_),
    .Y(_10330_));
 sky130_fd_sc_hd__and3_1 _14605_ (.A(_10071_),
    .B(\line_cache[128][0] ),
    .C(_09758_),
    .X(_10331_));
 sky130_fd_sc_hd__a21o_1 _14606_ (.A1(\line_cache[129][0] ),
    .A2(_10330_),
    .B1(_10331_),
    .X(_10332_));
 sky130_fd_sc_hd__a221o_1 _14607_ (.A1(\line_cache[131][0] ),
    .A2(_10328_),
    .B1(\line_cache[130][0] ),
    .B2(_10329_),
    .C1(_10332_),
    .X(_10333_));
 sky130_fd_sc_hd__nor2_4 _14608_ (.A(_09760_),
    .B(_10268_),
    .Y(_10334_));
 sky130_fd_sc_hd__nor2_4 _14609_ (.A(_09760_),
    .B(_10115_),
    .Y(_10335_));
 sky130_fd_sc_hd__nor2_4 _14610_ (.A(_10040_),
    .B(_09760_),
    .Y(_10336_));
 sky130_fd_sc_hd__nor2_2 _14611_ (.A(_10032_),
    .B(_09760_),
    .Y(_10337_));
 sky130_fd_sc_hd__a22o_1 _14612_ (.A1(_10336_),
    .A2(\line_cache[140][0] ),
    .B1(\line_cache[141][0] ),
    .B2(_10337_),
    .X(_10338_));
 sky130_fd_sc_hd__a221o_1 _14613_ (.A1(\line_cache[143][0] ),
    .A2(_10334_),
    .B1(\line_cache[142][0] ),
    .B2(_10335_),
    .C1(_10338_),
    .X(_10339_));
 sky130_fd_sc_hd__nor2_2 _14614_ (.A(_10058_),
    .B(_09760_),
    .Y(_10340_));
 sky130_fd_sc_hd__nor2_2 _14615_ (.A(_09578_),
    .B(_09760_),
    .Y(_10341_));
 sky130_fd_sc_hd__nor2_2 _14616_ (.A(_10119_),
    .B(_09760_),
    .Y(_10342_));
 sky130_fd_sc_hd__nor2_2 _14617_ (.A(_09760_),
    .B(_10055_),
    .Y(_10343_));
 sky130_fd_sc_hd__a22o_1 _14618_ (.A1(_10342_),
    .A2(\line_cache[139][0] ),
    .B1(\line_cache[138][0] ),
    .B2(_10343_),
    .X(_10344_));
 sky130_fd_sc_hd__a221o_1 _14619_ (.A1(\line_cache[137][0] ),
    .A2(_10340_),
    .B1(\line_cache[136][0] ),
    .B2(_10341_),
    .C1(_10344_),
    .X(_10345_));
 sky130_fd_sc_hd__or4_1 _14620_ (.A(_10327_),
    .B(_10333_),
    .C(_10339_),
    .D(_10345_),
    .X(_10346_));
 sky130_fd_sc_hd__nor2_1 _14621_ (.A(_10321_),
    .B(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__nor2_4 _14622_ (.A(_09765_),
    .B(_10073_),
    .Y(_10348_));
 sky130_fd_sc_hd__nor2_2 _14623_ (.A(_09765_),
    .B(_10048_),
    .Y(_10349_));
 sky130_fd_sc_hd__and2_1 _14624_ (.A(_10349_),
    .B(\line_cache[99][0] ),
    .X(_10350_));
 sky130_fd_sc_hd__nor2_2 _14625_ (.A(_09765_),
    .B(_10069_),
    .Y(_10351_));
 sky130_fd_sc_hd__nor2_4 _14626_ (.A(_09765_),
    .B(_09569_),
    .Y(_10352_));
 sky130_fd_sc_hd__a22o_1 _14627_ (.A1(_10351_),
    .A2(\line_cache[96][0] ),
    .B1(_10352_),
    .B2(\line_cache[97][0] ),
    .X(_10353_));
 sky130_fd_sc_hd__a211o_1 _14628_ (.A1(\line_cache[98][0] ),
    .A2(_10348_),
    .B1(_10350_),
    .C1(_10353_),
    .X(_10354_));
 sky130_fd_sc_hd__inv_2 _14629_ (.A(_09765_),
    .Y(_10355_));
 sky130_fd_sc_hd__buf_4 _14630_ (.A(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__and3_1 _14631_ (.A(_10035_),
    .B(\line_cache[107][0] ),
    .C(_10356_),
    .X(_10357_));
 sky130_fd_sc_hd__and3_1 _14632_ (.A(_10176_),
    .B(\line_cache[105][0] ),
    .C(_10356_),
    .X(_10358_));
 sky130_fd_sc_hd__and3_1 _14633_ (.A(_10054_),
    .B(\line_cache[106][0] ),
    .C(_10356_),
    .X(_10359_));
 sky130_fd_sc_hd__inv_2 _14634_ (.A(_09578_),
    .Y(_10360_));
 sky130_fd_sc_hd__and3_1 _14635_ (.A(_10360_),
    .B(\line_cache[104][0] ),
    .C(_10356_),
    .X(_10361_));
 sky130_fd_sc_hd__or4_1 _14636_ (.A(_10357_),
    .B(_10358_),
    .C(_10359_),
    .D(_10361_),
    .X(_10362_));
 sky130_fd_sc_hd__and3_4 _14637_ (.A(_10356_),
    .B(_09531_),
    .C(_10109_),
    .X(_10363_));
 sky130_fd_sc_hd__nor2_4 _14638_ (.A(_09765_),
    .B(_10115_),
    .Y(_10364_));
 sky130_fd_sc_hd__nor2_4 _14639_ (.A(_09765_),
    .B(_10040_),
    .Y(_10365_));
 sky130_fd_sc_hd__nor2_4 _14640_ (.A(_09765_),
    .B(_10032_),
    .Y(_10366_));
 sky130_fd_sc_hd__a22o_1 _14641_ (.A1(_10365_),
    .A2(\line_cache[108][0] ),
    .B1(_10366_),
    .B2(\line_cache[109][0] ),
    .X(_10367_));
 sky130_fd_sc_hd__a221o_1 _14642_ (.A1(\line_cache[111][0] ),
    .A2(_10363_),
    .B1(\line_cache[110][0] ),
    .B2(_10364_),
    .C1(_10367_),
    .X(_10368_));
 sky130_fd_sc_hd__nor2_4 _14643_ (.A(_09765_),
    .B(_10062_),
    .Y(_10369_));
 sky130_fd_sc_hd__nor2_4 _14644_ (.A(_09765_),
    .B(_10045_),
    .Y(_10370_));
 sky130_fd_sc_hd__nor2_2 _14645_ (.A(_09765_),
    .B(_10050_),
    .Y(_10371_));
 sky130_fd_sc_hd__nor2_4 _14646_ (.A(_09765_),
    .B(_09596_),
    .Y(_10372_));
 sky130_fd_sc_hd__a22o_1 _14647_ (.A1(_10371_),
    .A2(\line_cache[100][0] ),
    .B1(_10372_),
    .B2(\line_cache[101][0] ),
    .X(_10373_));
 sky130_fd_sc_hd__a221o_1 _14648_ (.A1(\line_cache[103][0] ),
    .A2(_10369_),
    .B1(\line_cache[102][0] ),
    .B2(_10370_),
    .C1(_10373_),
    .X(_10374_));
 sky130_fd_sc_hd__or4_1 _14649_ (.A(_10354_),
    .B(_10362_),
    .C(_10368_),
    .D(_10374_),
    .X(_10375_));
 sky130_fd_sc_hd__nor2_4 _14650_ (.A(_09764_),
    .B(_10048_),
    .Y(_10376_));
 sky130_fd_sc_hd__nor2_4 _14651_ (.A(_09764_),
    .B(_10073_),
    .Y(_10377_));
 sky130_fd_sc_hd__nor2_2 _14652_ (.A(_09764_),
    .B(_10069_),
    .Y(_10378_));
 sky130_fd_sc_hd__nor2_2 _14653_ (.A(_09764_),
    .B(_09569_),
    .Y(_10379_));
 sky130_fd_sc_hd__a22o_1 _14654_ (.A1(_10378_),
    .A2(\line_cache[80][0] ),
    .B1(_10379_),
    .B2(\line_cache[81][0] ),
    .X(_10380_));
 sky130_fd_sc_hd__a221o_1 _14655_ (.A1(\line_cache[83][0] ),
    .A2(_10376_),
    .B1(\line_cache[82][0] ),
    .B2(_10377_),
    .C1(_10380_),
    .X(_10381_));
 sky130_fd_sc_hd__nor3_2 _14656_ (.A(_09546_),
    .B(_09764_),
    .C(_09601_),
    .Y(_10382_));
 sky130_fd_sc_hd__nor2_4 _14657_ (.A(_09764_),
    .B(_10115_),
    .Y(_10383_));
 sky130_fd_sc_hd__nor2_4 _14658_ (.A(_09764_),
    .B(_10040_),
    .Y(_10384_));
 sky130_fd_sc_hd__nor2_4 _14659_ (.A(_09764_),
    .B(_10032_),
    .Y(_10385_));
 sky130_fd_sc_hd__a22o_1 _14660_ (.A1(_10384_),
    .A2(\line_cache[92][0] ),
    .B1(_10385_),
    .B2(\line_cache[93][0] ),
    .X(_10386_));
 sky130_fd_sc_hd__a221o_1 _14661_ (.A1(\line_cache[95][0] ),
    .A2(net136),
    .B1(\line_cache[94][0] ),
    .B2(_10383_),
    .C1(_10386_),
    .X(_10387_));
 sky130_fd_sc_hd__nor2_2 _14662_ (.A(_09764_),
    .B(_10062_),
    .Y(_10388_));
 sky130_fd_sc_hd__nor2_4 _14663_ (.A(_09764_),
    .B(_10045_),
    .Y(_10389_));
 sky130_fd_sc_hd__nor2_4 _14664_ (.A(_09763_),
    .B(_10050_),
    .Y(_10390_));
 sky130_fd_sc_hd__nor2_4 _14665_ (.A(_09764_),
    .B(_09596_),
    .Y(_10391_));
 sky130_fd_sc_hd__a22o_1 _14666_ (.A1(_10390_),
    .A2(\line_cache[84][0] ),
    .B1(_10391_),
    .B2(\line_cache[85][0] ),
    .X(_10392_));
 sky130_fd_sc_hd__a221o_1 _14667_ (.A1(\line_cache[87][0] ),
    .A2(_10388_),
    .B1(\line_cache[86][0] ),
    .B2(_10389_),
    .C1(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__nor2_4 _14668_ (.A(_09764_),
    .B(_10119_),
    .Y(_10394_));
 sky130_fd_sc_hd__nor2_4 _14669_ (.A(_09764_),
    .B(_10055_),
    .Y(_10395_));
 sky130_fd_sc_hd__nor2_4 _14670_ (.A(_09764_),
    .B(_09578_),
    .Y(_10396_));
 sky130_fd_sc_hd__nor2_4 _14671_ (.A(_09764_),
    .B(_10058_),
    .Y(_10397_));
 sky130_fd_sc_hd__a22o_1 _14672_ (.A1(_10396_),
    .A2(\line_cache[88][0] ),
    .B1(_10397_),
    .B2(\line_cache[89][0] ),
    .X(_10398_));
 sky130_fd_sc_hd__a221o_1 _14673_ (.A1(\line_cache[91][0] ),
    .A2(_10394_),
    .B1(\line_cache[90][0] ),
    .B2(_10395_),
    .C1(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__or4_1 _14674_ (.A(_10381_),
    .B(_10387_),
    .C(_10393_),
    .D(_10399_),
    .X(_10400_));
 sky130_fd_sc_hd__nor2_1 _14675_ (.A(_10375_),
    .B(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__and3_2 _14676_ (.A(_10295_),
    .B(_10347_),
    .C(_10401_),
    .X(_10402_));
 sky130_fd_sc_hd__nand3_1 _14677_ (.A(_09986_),
    .B(_10216_),
    .C(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__a21oi_1 _14678_ (.A1(\line_cache[0][0] ),
    .A2(_09912_),
    .B1(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__nor2_4 _14679_ (.A(_08979_),
    .B(_10404_),
    .Y(net126));
 sky130_fd_sc_hd__and2_1 _14680_ (.A(_09912_),
    .B(\line_cache[0][1] ),
    .X(_10405_));
 sky130_fd_sc_hd__and3_1 _14681_ (.A(_10102_),
    .B(\line_cache[70][1] ),
    .C(_10161_),
    .X(_10406_));
 sky130_fd_sc_hd__a22o_1 _14682_ (.A1(_10163_),
    .A2(\line_cache[68][1] ),
    .B1(_10164_),
    .B2(\line_cache[69][1] ),
    .X(_10407_));
 sky130_fd_sc_hd__a211o_1 _14683_ (.A1(\line_cache[71][1] ),
    .A2(_10159_),
    .B1(_10406_),
    .C1(_10407_),
    .X(_10408_));
 sky130_fd_sc_hd__and3_1 _14684_ (.A(_10031_),
    .B(\line_cache[77][1] ),
    .C(_10167_),
    .X(_10409_));
 sky130_fd_sc_hd__and3_1 _14685_ (.A(_10038_),
    .B(\line_cache[78][1] ),
    .C(_10167_),
    .X(_10410_));
 sky130_fd_sc_hd__and3_1 _14686_ (.A(_10041_),
    .B(\line_cache[76][1] ),
    .C(_10161_),
    .X(_10411_));
 sky130_fd_sc_hd__a2111o_1 _14687_ (.A1(_10168_),
    .A2(\line_cache[79][1] ),
    .B1(_10409_),
    .C1(_10410_),
    .D1(_10411_),
    .X(_10412_));
 sky130_fd_sc_hd__and3_1 _14688_ (.A(_10176_),
    .B(\line_cache[73][1] ),
    .C(_10167_),
    .X(_10413_));
 sky130_fd_sc_hd__a21o_1 _14689_ (.A1(\line_cache[72][1] ),
    .A2(_10175_),
    .B1(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__a221o_1 _14690_ (.A1(\line_cache[75][1] ),
    .A2(_10173_),
    .B1(\line_cache[74][1] ),
    .B2(_10174_),
    .C1(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__a22o_1 _14691_ (.A1(_10182_),
    .A2(\line_cache[64][1] ),
    .B1(_10183_),
    .B2(\line_cache[65][1] ),
    .X(_10416_));
 sky130_fd_sc_hd__a221o_1 _14692_ (.A1(\line_cache[67][1] ),
    .A2(_10180_),
    .B1(\line_cache[66][1] ),
    .B2(_10181_),
    .C1(_10416_),
    .X(_10417_));
 sky130_fd_sc_hd__or4_2 _14693_ (.A(_10408_),
    .B(_10412_),
    .C(_10415_),
    .D(_10417_),
    .X(_10418_));
 sky130_fd_sc_hd__a22o_1 _14694_ (.A1(_10189_),
    .A2(\line_cache[252][1] ),
    .B1(_10190_),
    .B2(\line_cache[251][1] ),
    .X(_10419_));
 sky130_fd_sc_hd__a221o_1 _14695_ (.A1(\line_cache[254][1] ),
    .A2(_10187_),
    .B1(\line_cache[253][1] ),
    .B2(_10188_),
    .C1(_10419_),
    .X(_10420_));
 sky130_fd_sc_hd__a22o_1 _14696_ (.A1(_10195_),
    .A2(\line_cache[248][1] ),
    .B1(_10196_),
    .B2(\line_cache[247][1] ),
    .X(_10421_));
 sky130_fd_sc_hd__a221o_1 _14697_ (.A1(\line_cache[250][1] ),
    .A2(_10193_),
    .B1(\line_cache[249][1] ),
    .B2(_10194_),
    .C1(_10421_),
    .X(_10422_));
 sky130_fd_sc_hd__and2b_1 _14698_ (.A_N(_10200_),
    .B(\line_cache[240][1] ),
    .X(_10423_));
 sky130_fd_sc_hd__and2b_1 _14699_ (.A_N(_09570_),
    .B(\line_cache[241][1] ),
    .X(_10424_));
 sky130_fd_sc_hd__and2b_1 _14700_ (.A_N(_10203_),
    .B(\line_cache[242][1] ),
    .X(_10425_));
 sky130_fd_sc_hd__a2111o_1 _14701_ (.A1(\line_cache[239][1] ),
    .A2(_10199_),
    .B1(_10423_),
    .C1(_10424_),
    .D1(_10425_),
    .X(_10426_));
 sky130_fd_sc_hd__and2b_1 _14702_ (.A_N(_10206_),
    .B(\line_cache[243][1] ),
    .X(_10427_));
 sky130_fd_sc_hd__and2b_1 _14703_ (.A_N(_10208_),
    .B(\line_cache[244][1] ),
    .X(_10428_));
 sky130_fd_sc_hd__and2b_1 _14704_ (.A_N(_09597_),
    .B(\line_cache[245][1] ),
    .X(_10429_));
 sky130_fd_sc_hd__and2b_1 _14705_ (.A_N(_10211_),
    .B(\line_cache[246][1] ),
    .X(_10430_));
 sky130_fd_sc_hd__or4_1 _14706_ (.A(_10427_),
    .B(_10428_),
    .C(_10429_),
    .D(_10430_),
    .X(_10431_));
 sky130_fd_sc_hd__or4_1 _14707_ (.A(_10420_),
    .B(_10422_),
    .C(_10426_),
    .D(_10431_),
    .X(_10432_));
 sky130_fd_sc_hd__and3_1 _14708_ (.A(_09595_),
    .B(\line_cache[229][1] ),
    .C(_10099_),
    .X(_10433_));
 sky130_fd_sc_hd__clkbuf_4 _14709_ (.A(_10099_),
    .X(_10434_));
 sky130_fd_sc_hd__and3_1 _14710_ (.A(_10102_),
    .B(\line_cache[230][1] ),
    .C(_10434_),
    .X(_10435_));
 sky130_fd_sc_hd__and3_1 _14711_ (.A(_10104_),
    .B(\line_cache[227][1] ),
    .C(_10434_),
    .X(_10436_));
 sky130_fd_sc_hd__clkbuf_4 _14712_ (.A(_10099_),
    .X(_10437_));
 sky130_fd_sc_hd__and3_1 _14713_ (.A(_10106_),
    .B(\line_cache[228][1] ),
    .C(_10437_),
    .X(_10438_));
 sky130_fd_sc_hd__or4_1 _14714_ (.A(_10433_),
    .B(_10435_),
    .C(_10436_),
    .D(_10438_),
    .X(_10439_));
 sky130_fd_sc_hd__and3_1 _14715_ (.A(_09544_),
    .B(\line_cache[223][1] ),
    .C(_10109_),
    .X(_10440_));
 sky130_fd_sc_hd__and3_1 _14716_ (.A(_10071_),
    .B(\line_cache[224][1] ),
    .C(_10434_),
    .X(_10441_));
 sky130_fd_sc_hd__and3_1 _14717_ (.A(_10067_),
    .B(\line_cache[225][1] ),
    .C(_10437_),
    .X(_10442_));
 sky130_fd_sc_hd__and3_1 _14718_ (.A(_10074_),
    .B(\line_cache[226][1] ),
    .C(_10100_),
    .X(_10443_));
 sky130_fd_sc_hd__or4_1 _14719_ (.A(_10440_),
    .B(_10441_),
    .C(_10442_),
    .D(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__a22o_1 _14720_ (.A1(_10118_),
    .A2(\line_cache[236][1] ),
    .B1(_10120_),
    .B2(\line_cache[235][1] ),
    .X(_10445_));
 sky130_fd_sc_hd__a221o_1 _14721_ (.A1(\line_cache[238][1] ),
    .A2(_10116_),
    .B1(\line_cache[237][1] ),
    .B2(_10117_),
    .C1(_10445_),
    .X(_10446_));
 sky130_fd_sc_hd__a22o_1 _14722_ (.A1(_10125_),
    .A2(\line_cache[232][1] ),
    .B1(_10126_),
    .B2(\line_cache[231][1] ),
    .X(_10447_));
 sky130_fd_sc_hd__a221o_1 _14723_ (.A1(\line_cache[234][1] ),
    .A2(_10123_),
    .B1(\line_cache[233][1] ),
    .B2(_10124_),
    .C1(_10447_),
    .X(_10448_));
 sky130_fd_sc_hd__or4_1 _14724_ (.A(_10439_),
    .B(_10444_),
    .C(_10446_),
    .D(_10448_),
    .X(_10449_));
 sky130_fd_sc_hd__a22o_1 _14725_ (.A1(_10132_),
    .A2(\line_cache[220][1] ),
    .B1(_10133_),
    .B2(\line_cache[219][1] ),
    .X(_10450_));
 sky130_fd_sc_hd__a221o_1 _14726_ (.A1(\line_cache[222][1] ),
    .A2(_10130_),
    .B1(\line_cache[221][1] ),
    .B2(_10131_),
    .C1(_10450_),
    .X(_10451_));
 sky130_fd_sc_hd__a22o_1 _14727_ (.A1(_10138_),
    .A2(\line_cache[208][1] ),
    .B1(_10139_),
    .B2(\line_cache[207][1] ),
    .X(_10452_));
 sky130_fd_sc_hd__a221o_1 _14728_ (.A1(\line_cache[210][1] ),
    .A2(_10136_),
    .B1(\line_cache[209][1] ),
    .B2(_10137_),
    .C1(_10452_),
    .X(_10453_));
 sky130_fd_sc_hd__a22o_1 _14729_ (.A1(_10144_),
    .A2(\line_cache[216][1] ),
    .B1(_10145_),
    .B2(\line_cache[215][1] ),
    .X(_10454_));
 sky130_fd_sc_hd__a221o_1 _14730_ (.A1(\line_cache[218][1] ),
    .A2(_10142_),
    .B1(\line_cache[217][1] ),
    .B2(_10143_),
    .C1(_10454_),
    .X(_10455_));
 sky130_fd_sc_hd__and2b_1 _14731_ (.A_N(_10148_),
    .B(\line_cache[211][1] ),
    .X(_10456_));
 sky130_fd_sc_hd__nor2b_1 _14732_ (.A(_10150_),
    .B_N(\line_cache[212][1] ),
    .Y(_10457_));
 sky130_fd_sc_hd__and2b_1 _14733_ (.A_N(_10152_),
    .B(\line_cache[213][1] ),
    .X(_10458_));
 sky130_fd_sc_hd__and2b_1 _14734_ (.A_N(_10154_),
    .B(\line_cache[214][1] ),
    .X(_10459_));
 sky130_fd_sc_hd__or4_1 _14735_ (.A(_10456_),
    .B(_10457_),
    .C(_10458_),
    .D(_10459_),
    .X(_10460_));
 sky130_fd_sc_hd__or4_1 _14736_ (.A(_10451_),
    .B(_10453_),
    .C(_10455_),
    .D(_10460_),
    .X(_10461_));
 sky130_fd_sc_hd__or2_1 _14737_ (.A(_10449_),
    .B(_10461_),
    .X(_10462_));
 sky130_fd_sc_hd__or3_2 _14738_ (.A(_10418_),
    .B(_10432_),
    .C(_10462_),
    .X(_10463_));
 sky130_fd_sc_hd__and3_1 _14739_ (.A(_10035_),
    .B(\line_cache[203][1] ),
    .C(_09539_),
    .X(_10464_));
 sky130_fd_sc_hd__and3_1 _14740_ (.A(_10038_),
    .B(\line_cache[206][1] ),
    .C(_10075_),
    .X(_10465_));
 sky130_fd_sc_hd__and3_1 _14741_ (.A(_10041_),
    .B(\line_cache[204][1] ),
    .C(_10075_),
    .X(_10466_));
 sky130_fd_sc_hd__a2111o_1 _14742_ (.A1(\line_cache[205][1] ),
    .A2(_10033_),
    .B1(_10464_),
    .C1(_10465_),
    .D1(_10466_),
    .X(_10467_));
 sky130_fd_sc_hd__a22o_1 _14743_ (.A1(_10049_),
    .A2(\line_cache[195][1] ),
    .B1(\line_cache[196][1] ),
    .B2(_10051_),
    .X(_10468_));
 sky130_fd_sc_hd__a221o_1 _14744_ (.A1(\line_cache[198][1] ),
    .A2(_10046_),
    .B1(\line_cache[197][1] ),
    .B2(_10047_),
    .C1(_10468_),
    .X(_10469_));
 sky130_fd_sc_hd__a22o_1 _14745_ (.A1(_10060_),
    .A2(\line_cache[200][1] ),
    .B1(_10063_),
    .B2(\line_cache[199][1] ),
    .X(_10470_));
 sky130_fd_sc_hd__a221o_1 _14746_ (.A1(\line_cache[202][1] ),
    .A2(_10056_),
    .B1(\line_cache[201][1] ),
    .B2(_10059_),
    .C1(_10470_),
    .X(_10471_));
 sky130_fd_sc_hd__and3_1 _14747_ (.A(_10067_),
    .B(\line_cache[193][1] ),
    .C(_09540_),
    .X(_10472_));
 sky130_fd_sc_hd__and3_1 _14748_ (.A(_10071_),
    .B(\line_cache[192][1] ),
    .C(_09540_),
    .X(_10473_));
 sky130_fd_sc_hd__and3_1 _14749_ (.A(_10074_),
    .B(\line_cache[194][1] ),
    .C(_09540_),
    .X(_10474_));
 sky130_fd_sc_hd__a2111o_1 _14750_ (.A1(_10066_),
    .A2(\line_cache[286][1] ),
    .B1(_10472_),
    .C1(_10473_),
    .D1(_10474_),
    .X(_10475_));
 sky130_fd_sc_hd__or4_1 _14751_ (.A(_10467_),
    .B(_10469_),
    .C(_10471_),
    .D(_10475_),
    .X(_10476_));
 sky130_fd_sc_hd__a22o_1 _14752_ (.A1(_09623_),
    .A2(\line_cache[275][1] ),
    .B1(_09620_),
    .B2(\line_cache[274][1] ),
    .X(_10477_));
 sky130_fd_sc_hd__a22o_1 _14753_ (.A1(_10080_),
    .A2(\line_cache[276][1] ),
    .B1(\line_cache[277][1] ),
    .B2(_10081_),
    .X(_10478_));
 sky130_fd_sc_hd__a22o_1 _14754_ (.A1(_10086_),
    .A2(\line_cache[270][1] ),
    .B1(\line_cache[269][1] ),
    .B2(_10088_),
    .X(_10479_));
 sky130_fd_sc_hd__a221o_1 _14755_ (.A1(\line_cache[273][1] ),
    .A2(_10083_),
    .B1(\line_cache[272][1] ),
    .B2(_10084_),
    .C1(_10479_),
    .X(_10480_));
 sky130_fd_sc_hd__a22o_1 _14756_ (.A1(_09658_),
    .A2(\line_cache[283][1] ),
    .B1(\line_cache[282][1] ),
    .B2(_09661_),
    .X(_10481_));
 sky130_fd_sc_hd__a22o_1 _14757_ (.A1(_09645_),
    .A2(\line_cache[285][1] ),
    .B1(\line_cache[284][1] ),
    .B2(_09648_),
    .X(_10482_));
 sky130_fd_sc_hd__a22o_1 _14758_ (.A1(_09639_),
    .A2(\line_cache[279][1] ),
    .B1(\line_cache[278][1] ),
    .B2(_09636_),
    .X(_10483_));
 sky130_fd_sc_hd__a221o_1 _14759_ (.A1(\line_cache[281][1] ),
    .A2(_09663_),
    .B1(\line_cache[280][1] ),
    .B2(_09655_),
    .C1(_10483_),
    .X(_10484_));
 sky130_fd_sc_hd__or3_1 _14760_ (.A(_10481_),
    .B(_10482_),
    .C(_10484_),
    .X(_10485_));
 sky130_fd_sc_hd__or4_1 _14761_ (.A(_10477_),
    .B(_10478_),
    .C(_10480_),
    .D(_10485_),
    .X(_10486_));
 sky130_fd_sc_hd__nor2_1 _14762_ (.A(_10476_),
    .B(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__and2b_1 _14763_ (.A_N(_09987_),
    .B(\line_cache[256][1] ),
    .X(_10488_));
 sky130_fd_sc_hd__and2b_1 _14764_ (.A_N(_09747_),
    .B(\line_cache[302][1] ),
    .X(_10489_));
 sky130_fd_sc_hd__a22o_1 _14765_ (.A1(_09743_),
    .A2(\line_cache[301][1] ),
    .B1(\line_cache[300][1] ),
    .B2(_09742_),
    .X(_10490_));
 sky130_fd_sc_hd__or3_1 _14766_ (.A(_10488_),
    .B(_10489_),
    .C(_10490_),
    .X(_10491_));
 sky130_fd_sc_hd__and3_1 _14767_ (.A(_09917_),
    .B(_09691_),
    .C(\line_cache[258][1] ),
    .X(_10492_));
 sky130_fd_sc_hd__and3_1 _14768_ (.A(_09848_),
    .B(_09691_),
    .C(\line_cache[260][1] ),
    .X(_10493_));
 sky130_fd_sc_hd__and3_1 _14769_ (.A(_09919_),
    .B(_09611_),
    .C(\line_cache[257][1] ),
    .X(_10494_));
 sky130_fd_sc_hd__and3_1 _14770_ (.A(_09840_),
    .B(_09611_),
    .C(\line_cache[259][1] ),
    .X(_10495_));
 sky130_fd_sc_hd__or4_1 _14771_ (.A(_10492_),
    .B(_10493_),
    .C(_10494_),
    .D(_10495_),
    .X(_10496_));
 sky130_fd_sc_hd__and3_1 _14772_ (.A(_09858_),
    .B(_09547_),
    .C(\line_cache[267][1] ),
    .X(_10497_));
 sky130_fd_sc_hd__a22o_1 _14773_ (.A1(_09998_),
    .A2(\line_cache[265][1] ),
    .B1(\line_cache[266][1] ),
    .B2(_09999_),
    .X(_10498_));
 sky130_fd_sc_hd__a311o_1 _14774_ (.A1(_09548_),
    .A2(\line_cache[268][1] ),
    .A3(_09862_),
    .B1(_10497_),
    .C1(_10498_),
    .X(_10499_));
 sky130_fd_sc_hd__nand2_1 _14775_ (.A(_10007_),
    .B(\line_cache[262][1] ),
    .Y(_10500_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(_10010_),
    .B(\line_cache[261][1] ),
    .Y(_10501_));
 sky130_fd_sc_hd__nand2_1 _14777_ (.A(_10500_),
    .B(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__a221oi_1 _14778_ (.A1(_10003_),
    .A2(\line_cache[264][1] ),
    .B1(_10005_),
    .B2(\line_cache[263][1] ),
    .C1(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__or4b_1 _14779_ (.A(_10491_),
    .B(_10496_),
    .C(_10499_),
    .D_N(_10503_),
    .X(_10504_));
 sky130_fd_sc_hd__a22o_1 _14780_ (.A1(_09682_),
    .A2(\line_cache[308][1] ),
    .B1(\line_cache[309][1] ),
    .B2(_09685_),
    .X(_10505_));
 sky130_fd_sc_hd__a221o_1 _14781_ (.A1(\line_cache[311][1] ),
    .A2(_09689_),
    .B1(\line_cache[310][1] ),
    .B2(_09693_),
    .C1(_10505_),
    .X(_10506_));
 sky130_fd_sc_hd__a22o_1 _14782_ (.A1(_09728_),
    .A2(\line_cache[295][1] ),
    .B1(\line_cache[294][1] ),
    .B2(_09726_),
    .X(_10507_));
 sky130_fd_sc_hd__a221o_1 _14783_ (.A1(\line_cache[293][1] ),
    .A2(_09730_),
    .B1(\line_cache[292][1] ),
    .B2(_10018_),
    .C1(_10507_),
    .X(_10508_));
 sky130_fd_sc_hd__a22o_1 _14784_ (.A1(_09716_),
    .A2(\line_cache[296][1] ),
    .B1(\line_cache[297][1] ),
    .B2(_09721_),
    .X(_10509_));
 sky130_fd_sc_hd__a221o_1 _14785_ (.A1(\line_cache[299][1] ),
    .A2(_09718_),
    .B1(\line_cache[298][1] ),
    .B2(_09720_),
    .C1(_10509_),
    .X(_10510_));
 sky130_fd_sc_hd__a22o_1 _14786_ (.A1(_10025_),
    .A2(\line_cache[288][1] ),
    .B1(\line_cache[289][1] ),
    .B2(_10026_),
    .X(_10511_));
 sky130_fd_sc_hd__a221o_1 _14787_ (.A1(\line_cache[291][1] ),
    .A2(_10023_),
    .B1(\line_cache[290][1] ),
    .B2(_10024_),
    .C1(_10511_),
    .X(_10512_));
 sky130_fd_sc_hd__or4_2 _14788_ (.A(_10506_),
    .B(_10508_),
    .C(_10510_),
    .D(_10512_),
    .X(_10513_));
 sky130_fd_sc_hd__nor2_1 _14789_ (.A(_10504_),
    .B(_10513_),
    .Y(_10514_));
 sky130_fd_sc_hd__nand2_1 _14790_ (.A(_10487_),
    .B(_10514_),
    .Y(_10515_));
 sky130_fd_sc_hd__nor2_1 _14791_ (.A(_10463_),
    .B(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__a22o_1 _14792_ (.A1(_09842_),
    .A2(\line_cache[6][1] ),
    .B1(\line_cache[5][1] ),
    .B2(_09844_),
    .X(_10517_));
 sky130_fd_sc_hd__a221o_1 _14793_ (.A1(\line_cache[4][1] ),
    .A2(_09850_),
    .B1(\line_cache[3][1] ),
    .B2(_09914_),
    .C1(_10517_),
    .X(_10518_));
 sky130_fd_sc_hd__and3_1 _14794_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][1] ),
    .X(_10519_));
 sky130_fd_sc_hd__and3_1 _14795_ (.A(_09919_),
    .B(_09533_),
    .C(\line_cache[1][1] ),
    .X(_10520_));
 sky130_fd_sc_hd__a211o_1 _14796_ (.A1(\line_cache[15][1] ),
    .A2(_09867_),
    .B1(_10519_),
    .C1(_10520_),
    .X(_10521_));
 sky130_fd_sc_hd__and3_1 _14797_ (.A(_09922_),
    .B(_09532_),
    .C(\line_cache[63][1] ),
    .X(_10522_));
 sky130_fd_sc_hd__a31o_1 _14798_ (.A1(_09548_),
    .A2(\line_cache[319][1] ),
    .A3(_09922_),
    .B1(_10522_),
    .X(_10523_));
 sky130_fd_sc_hd__a221o_1 _14799_ (.A1(\line_cache[47][1] ),
    .A2(_09806_),
    .B1(\line_cache[31][1] ),
    .B2(_09907_),
    .C1(_10523_),
    .X(_10524_));
 sky130_fd_sc_hd__nand2_1 _14800_ (.A(_09746_),
    .B(\line_cache[303][1] ),
    .Y(_10525_));
 sky130_fd_sc_hd__nand2_1 _14801_ (.A(_09930_),
    .B(\line_cache[271][1] ),
    .Y(_10526_));
 sky130_fd_sc_hd__nand2_1 _14802_ (.A(_10525_),
    .B(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__a221oi_2 _14803_ (.A1(\line_cache[255][1] ),
    .A2(_09926_),
    .B1(\line_cache[287][1] ),
    .B2(_09927_),
    .C1(_10527_),
    .Y(_10528_));
 sky130_fd_sc_hd__or4b_1 _14804_ (.A(_10518_),
    .B(_10521_),
    .C(_10524_),
    .D_N(_10528_),
    .X(_10529_));
 sky130_fd_sc_hd__a22o_1 _14805_ (.A1(_09803_),
    .A2(\line_cache[45][1] ),
    .B1(\line_cache[46][1] ),
    .B2(_09804_),
    .X(_10530_));
 sky130_fd_sc_hd__a22o_1 _14806_ (.A1(_09824_),
    .A2(\line_cache[48][1] ),
    .B1(\line_cache[49][1] ),
    .B2(_09826_),
    .X(_10531_));
 sky130_fd_sc_hd__nand2_1 _14807_ (.A(_09787_),
    .B(\line_cache[41][1] ),
    .Y(_10532_));
 sky130_fd_sc_hd__nand2_1 _14808_ (.A(_09789_),
    .B(\line_cache[42][1] ),
    .Y(_10533_));
 sky130_fd_sc_hd__nand2_1 _14809_ (.A(_10532_),
    .B(_10533_),
    .Y(_10534_));
 sky130_fd_sc_hd__a221oi_2 _14810_ (.A1(_09785_),
    .A2(\line_cache[43][1] ),
    .B1(\line_cache[44][1] ),
    .B2(_09801_),
    .C1(_10534_),
    .Y(_10535_));
 sky130_fd_sc_hd__or3b_1 _14811_ (.A(_10530_),
    .B(_10531_),
    .C_N(_10535_),
    .X(_10536_));
 sky130_fd_sc_hd__a22o_1 _14812_ (.A1(_09699_),
    .A2(\line_cache[317][1] ),
    .B1(\line_cache[316][1] ),
    .B2(_09697_),
    .X(_10537_));
 sky130_fd_sc_hd__a22o_1 _14813_ (.A1(_09832_),
    .A2(\line_cache[58][1] ),
    .B1(\line_cache[59][1] ),
    .B2(_09833_),
    .X(_10538_));
 sky130_fd_sc_hd__a22o_1 _14814_ (.A1(_09819_),
    .A2(\line_cache[61][1] ),
    .B1(\line_cache[60][1] ),
    .B2(_09817_),
    .X(_10539_));
 sky130_fd_sc_hd__a22o_1 _14815_ (.A1(_09822_),
    .A2(\line_cache[62][1] ),
    .B1(\line_cache[318][1] ),
    .B2(_09702_),
    .X(_10540_));
 sky130_fd_sc_hd__or4_1 _14816_ (.A(_10537_),
    .B(_10538_),
    .C(_10539_),
    .D(_10540_),
    .X(_10541_));
 sky130_fd_sc_hd__a22o_1 _14817_ (.A1(_09675_),
    .A2(\line_cache[304][1] ),
    .B1(\line_cache[305][1] ),
    .B2(_09676_),
    .X(_10542_));
 sky130_fd_sc_hd__a22o_1 _14818_ (.A1(_09705_),
    .A2(\line_cache[312][1] ),
    .B1(\line_cache[313][1] ),
    .B2(_09707_),
    .X(_10543_));
 sky130_fd_sc_hd__a22o_1 _14819_ (.A1(_09708_),
    .A2(\line_cache[314][1] ),
    .B1(\line_cache[315][1] ),
    .B2(_09709_),
    .X(_10544_));
 sky130_fd_sc_hd__a22o_1 _14820_ (.A1(_09677_),
    .A2(\line_cache[306][1] ),
    .B1(\line_cache[307][1] ),
    .B2(_09678_),
    .X(_10545_));
 sky130_fd_sc_hd__or4_1 _14821_ (.A(_10542_),
    .B(_10543_),
    .C(_10544_),
    .D(_10545_),
    .X(_10546_));
 sky130_fd_sc_hd__a22o_1 _14822_ (.A1(_09830_),
    .A2(\line_cache[56][1] ),
    .B1(\line_cache[57][1] ),
    .B2(_09834_),
    .X(_10547_));
 sky130_fd_sc_hd__a22o_1 _14823_ (.A1(_09809_),
    .A2(\line_cache[52][1] ),
    .B1(\line_cache[53][1] ),
    .B2(_09811_),
    .X(_10548_));
 sky130_fd_sc_hd__a22o_1 _14824_ (.A1(_09827_),
    .A2(\line_cache[50][1] ),
    .B1(\line_cache[51][1] ),
    .B2(_09828_),
    .X(_10549_));
 sky130_fd_sc_hd__a22o_1 _14825_ (.A1(_09813_),
    .A2(\line_cache[54][1] ),
    .B1(\line_cache[55][1] ),
    .B2(_09815_),
    .X(_10550_));
 sky130_fd_sc_hd__or4_1 _14826_ (.A(_10547_),
    .B(_10548_),
    .C(_10549_),
    .D(_10550_),
    .X(_10551_));
 sky130_fd_sc_hd__or4_2 _14827_ (.A(_10536_),
    .B(_10541_),
    .C(_10546_),
    .D(_10551_),
    .X(_10552_));
 sky130_fd_sc_hd__nand2_1 _14828_ (.A(_09864_),
    .B(\line_cache[12][1] ),
    .Y(_10553_));
 sky130_fd_sc_hd__nand2_1 _14829_ (.A(_09860_),
    .B(\line_cache[11][1] ),
    .Y(_10554_));
 sky130_fd_sc_hd__nand2_1 _14830_ (.A(_10553_),
    .B(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__a221oi_2 _14831_ (.A1(_09870_),
    .A2(\line_cache[14][1] ),
    .B1(\line_cache[13][1] ),
    .B2(_09873_),
    .C1(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__nand2_1 _14832_ (.A(_09853_),
    .B(\line_cache[10][1] ),
    .Y(_10557_));
 sky130_fd_sc_hd__nand2_1 _14833_ (.A(_09857_),
    .B(\line_cache[9][1] ),
    .Y(_10558_));
 sky130_fd_sc_hd__nand2_1 _14834_ (.A(_10557_),
    .B(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__a221oi_1 _14835_ (.A1(_09855_),
    .A2(\line_cache[8][1] ),
    .B1(_09847_),
    .B2(\line_cache[7][1] ),
    .C1(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__nand2_1 _14836_ (.A(_10556_),
    .B(_10560_),
    .Y(_10561_));
 sky130_fd_sc_hd__and3_1 _14837_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][1] ),
    .X(_10562_));
 sky130_fd_sc_hd__a22o_1 _14838_ (.A1(_09884_),
    .A2(\line_cache[23][1] ),
    .B1(\line_cache[22][1] ),
    .B2(_09886_),
    .X(_10563_));
 sky130_fd_sc_hd__a22o_1 _14839_ (.A1(_09877_),
    .A2(\line_cache[19][1] ),
    .B1(\line_cache[18][1] ),
    .B2(_09878_),
    .X(_10564_));
 sky130_fd_sc_hd__a221o_1 _14840_ (.A1(\line_cache[17][1] ),
    .A2(_09969_),
    .B1(\line_cache[16][1] ),
    .B2(_09970_),
    .C1(_10564_),
    .X(_10565_));
 sky130_fd_sc_hd__a2111o_1 _14841_ (.A1(\line_cache[20][1] ),
    .A2(_09888_),
    .B1(_10562_),
    .C1(_10563_),
    .D1(_10565_),
    .X(_10566_));
 sky130_fd_sc_hd__a22o_1 _14842_ (.A1(_09796_),
    .A2(\line_cache[33][1] ),
    .B1(\line_cache[34][1] ),
    .B2(_09798_),
    .X(_10567_));
 sky130_fd_sc_hd__a221o_1 _14843_ (.A1(\line_cache[36][1] ),
    .A2(_09777_),
    .B1(\line_cache[35][1] ),
    .B2(_09794_),
    .C1(_10567_),
    .X(_10568_));
 sky130_fd_sc_hd__a22o_1 _14844_ (.A1(_09890_),
    .A2(\line_cache[27][1] ),
    .B1(\line_cache[26][1] ),
    .B2(_09896_),
    .X(_10569_));
 sky130_fd_sc_hd__a221oi_2 _14845_ (.A1(\line_cache[25][1] ),
    .A2(_09892_),
    .B1(\line_cache[24][1] ),
    .B2(_09895_),
    .C1(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__a22o_1 _14846_ (.A1(_09903_),
    .A2(\line_cache[29][1] ),
    .B1(\line_cache[28][1] ),
    .B2(_09900_),
    .X(_10571_));
 sky130_fd_sc_hd__a221oi_1 _14847_ (.A1(\line_cache[32][1] ),
    .A2(_09792_),
    .B1(\line_cache[30][1] ),
    .B2(_09905_),
    .C1(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__nand2_1 _14848_ (.A(_09773_),
    .B(\line_cache[38][1] ),
    .Y(_10573_));
 sky130_fd_sc_hd__nand2_1 _14849_ (.A(_09775_),
    .B(\line_cache[37][1] ),
    .Y(_10574_));
 sky130_fd_sc_hd__nand2_1 _14850_ (.A(_10573_),
    .B(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__a221oi_2 _14851_ (.A1(_09783_),
    .A2(\line_cache[40][1] ),
    .B1(\line_cache[39][1] ),
    .B2(_09780_),
    .C1(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__and4b_1 _14852_ (.A_N(_10568_),
    .B(_10570_),
    .C(_10572_),
    .D(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__or3b_2 _14853_ (.A(_10561_),
    .B(_10566_),
    .C_N(_10577_),
    .X(_10578_));
 sky130_fd_sc_hd__nor3_1 _14854_ (.A(_10529_),
    .B(_10552_),
    .C(_10578_),
    .Y(_10579_));
 sky130_fd_sc_hd__a22o_1 _14855_ (.A1(_10244_),
    .A2(\line_cache[173][1] ),
    .B1(\line_cache[172][1] ),
    .B2(_10245_),
    .X(_10580_));
 sky130_fd_sc_hd__a221o_1 _14856_ (.A1(\line_cache[175][1] ),
    .A2(_10242_),
    .B1(\line_cache[174][1] ),
    .B2(_10243_),
    .C1(_10580_),
    .X(_10581_));
 sky130_fd_sc_hd__a22o_1 _14857_ (.A1(_10263_),
    .A2(\line_cache[170][1] ),
    .B1(\line_cache[171][1] ),
    .B2(_10262_),
    .X(_10582_));
 sky130_fd_sc_hd__a221o_1 _14858_ (.A1(\line_cache[169][1] ),
    .A2(_10260_),
    .B1(\line_cache[168][1] ),
    .B2(_10261_),
    .C1(_10582_),
    .X(_10583_));
 sky130_fd_sc_hd__a22o_1 _14859_ (.A1(_10256_),
    .A2(\line_cache[160][1] ),
    .B1(\line_cache[161][1] ),
    .B2(_10257_),
    .X(_10584_));
 sky130_fd_sc_hd__and3_1 _14860_ (.A(_10104_),
    .B(_09751_),
    .C(\line_cache[163][1] ),
    .X(_10585_));
 sky130_fd_sc_hd__nand2_1 _14861_ (.A(_10249_),
    .B(\line_cache[166][1] ),
    .Y(_10586_));
 sky130_fd_sc_hd__nand2_1 _14862_ (.A(_10248_),
    .B(\line_cache[167][1] ),
    .Y(_10587_));
 sky130_fd_sc_hd__nand2_1 _14863_ (.A(_10586_),
    .B(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__a221o_1 _14864_ (.A1(\line_cache[165][1] ),
    .A2(_10250_),
    .B1(\line_cache[164][1] ),
    .B2(_10251_),
    .C1(_10588_),
    .X(_10589_));
 sky130_fd_sc_hd__a2111o_1 _14865_ (.A1(\line_cache[162][1] ),
    .A2(_10255_),
    .B1(_10584_),
    .C1(_10585_),
    .D1(_10589_),
    .X(_10590_));
 sky130_fd_sc_hd__nor3_1 _14866_ (.A(_10581_),
    .B(_10583_),
    .C(_10590_),
    .Y(_10591_));
 sky130_fd_sc_hd__a22o_1 _14867_ (.A1(_10275_),
    .A2(\line_cache[187][1] ),
    .B1(\line_cache[186][1] ),
    .B2(_10276_),
    .X(_10592_));
 sky130_fd_sc_hd__a221o_1 _14868_ (.A1(\line_cache[185][1] ),
    .A2(_10278_),
    .B1(\line_cache[184][1] ),
    .B2(_10277_),
    .C1(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__a22o_1 _14869_ (.A1(_10284_),
    .A2(\line_cache[176][1] ),
    .B1(_10285_),
    .B2(\line_cache[177][1] ),
    .X(_10594_));
 sky130_fd_sc_hd__a221oi_2 _14870_ (.A1(\line_cache[179][1] ),
    .A2(_10282_),
    .B1(\line_cache[178][1] ),
    .B2(_10283_),
    .C1(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__and3_1 _14871_ (.A(_10289_),
    .B(_10102_),
    .C(\line_cache[182][1] ),
    .X(_10596_));
 sky130_fd_sc_hd__and3_1 _14872_ (.A(_10288_),
    .B(_10098_),
    .C(\line_cache[181][1] ),
    .X(_10597_));
 sky130_fd_sc_hd__a31o_1 _14873_ (.A1(\line_cache[180][1] ),
    .A2(_10289_),
    .A3(_10106_),
    .B1(_10597_),
    .X(_10598_));
 sky130_fd_sc_hd__a311oi_1 _14874_ (.A1(\line_cache[183][1] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_10596_),
    .C1(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__a22o_1 _14875_ (.A1(_10272_),
    .A2(\line_cache[189][1] ),
    .B1(\line_cache[188][1] ),
    .B2(_10271_),
    .X(_10600_));
 sky130_fd_sc_hd__a221oi_1 _14876_ (.A1(\line_cache[191][1] ),
    .A2(_10269_),
    .B1(\line_cache[190][1] ),
    .B2(_10270_),
    .C1(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__and4b_1 _14877_ (.A_N(_10593_),
    .B(_10595_),
    .C(_10599_),
    .D(_10601_),
    .X(_10602_));
 sky130_fd_sc_hd__a22o_1 _14878_ (.A1(_10219_),
    .A2(\line_cache[157][1] ),
    .B1(\line_cache[156][1] ),
    .B2(_10220_),
    .X(_10603_));
 sky130_fd_sc_hd__a221o_1 _14879_ (.A1(\line_cache[159][1] ),
    .A2(_10217_),
    .B1(\line_cache[158][1] ),
    .B2(_10218_),
    .C1(_10603_),
    .X(_10604_));
 sky130_fd_sc_hd__a22o_1 _14880_ (.A1(_10238_),
    .A2(\line_cache[154][1] ),
    .B1(\line_cache[155][1] ),
    .B2(_10237_),
    .X(_10605_));
 sky130_fd_sc_hd__a221o_1 _14881_ (.A1(\line_cache[153][1] ),
    .A2(_10235_),
    .B1(\line_cache[152][1] ),
    .B2(_10236_),
    .C1(_10605_),
    .X(_10606_));
 sky130_fd_sc_hd__a22o_1 _14882_ (.A1(_10224_),
    .A2(\line_cache[148][1] ),
    .B1(\line_cache[149][1] ),
    .B2(_10223_),
    .X(_10607_));
 sky130_fd_sc_hd__a22o_1 _14883_ (.A1(_10225_),
    .A2(\line_cache[151][1] ),
    .B1(\line_cache[150][1] ),
    .B2(_10226_),
    .X(_10608_));
 sky130_fd_sc_hd__a22o_1 _14884_ (.A1(_10230_),
    .A2(\line_cache[144][1] ),
    .B1(\line_cache[145][1] ),
    .B2(_10229_),
    .X(_10609_));
 sky130_fd_sc_hd__a22o_1 _14885_ (.A1(_10231_),
    .A2(\line_cache[147][1] ),
    .B1(\line_cache[146][1] ),
    .B2(_10232_),
    .X(_10610_));
 sky130_fd_sc_hd__or4_1 _14886_ (.A(_10607_),
    .B(_10608_),
    .C(_10609_),
    .D(_10610_),
    .X(_10611_));
 sky130_fd_sc_hd__nor3_1 _14887_ (.A(_10604_),
    .B(_10606_),
    .C(_10611_),
    .Y(_10612_));
 sky130_fd_sc_hd__and3_2 _14888_ (.A(_10591_),
    .B(_10602_),
    .C(_10612_),
    .X(_10613_));
 sky130_fd_sc_hd__and3_1 _14889_ (.A(_10176_),
    .B(\line_cache[121][1] ),
    .C(_10302_),
    .X(_10614_));
 sky130_fd_sc_hd__a21o_1 _14890_ (.A1(\line_cache[120][1] ),
    .A2(_10317_),
    .B1(_10614_),
    .X(_10615_));
 sky130_fd_sc_hd__a221o_1 _14891_ (.A1(\line_cache[123][1] ),
    .A2(_10315_),
    .B1(\line_cache[122][1] ),
    .B2(_10316_),
    .C1(_10615_),
    .X(_10616_));
 sky130_fd_sc_hd__a22o_1 _14892_ (.A1(_10298_),
    .A2(\line_cache[112][1] ),
    .B1(_10299_),
    .B2(\line_cache[113][1] ),
    .X(_10617_));
 sky130_fd_sc_hd__a221o_1 _14893_ (.A1(\line_cache[115][1] ),
    .A2(_10296_),
    .B1(\line_cache[114][1] ),
    .B2(_10297_),
    .C1(_10617_),
    .X(_10618_));
 sky130_fd_sc_hd__a22o_1 _14894_ (.A1(_10311_),
    .A2(\line_cache[116][1] ),
    .B1(_10312_),
    .B2(\line_cache[117][1] ),
    .X(_10619_));
 sky130_fd_sc_hd__a221o_1 _14895_ (.A1(\line_cache[119][1] ),
    .A2(_10309_),
    .B1(\line_cache[118][1] ),
    .B2(_10310_),
    .C1(_10619_),
    .X(_10620_));
 sky130_fd_sc_hd__or3_2 _14896_ (.A(_09545_),
    .B(_09767_),
    .C(_09601_),
    .X(_10621_));
 sky130_fd_sc_hd__inv_2 _14897_ (.A(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__a22o_1 _14898_ (.A1(_10305_),
    .A2(\line_cache[124][1] ),
    .B1(_10306_),
    .B2(\line_cache[125][1] ),
    .X(_10623_));
 sky130_fd_sc_hd__a221o_1 _14899_ (.A1(\line_cache[126][1] ),
    .A2(_10304_),
    .B1(\line_cache[127][1] ),
    .B2(_10622_),
    .C1(_10623_),
    .X(_10624_));
 sky130_fd_sc_hd__or4_1 _14900_ (.A(_10616_),
    .B(_10618_),
    .C(_10620_),
    .D(_10624_),
    .X(_10625_));
 sky130_fd_sc_hd__nor2_1 _14901_ (.A(_09596_),
    .B(_09760_),
    .Y(_10626_));
 sky130_fd_sc_hd__a22o_1 _14902_ (.A1(_10322_),
    .A2(\line_cache[135][1] ),
    .B1(\line_cache[134][1] ),
    .B2(_10323_),
    .X(_10627_));
 sky130_fd_sc_hd__a221o_1 _14903_ (.A1(\line_cache[133][1] ),
    .A2(_10626_),
    .B1(\line_cache[132][1] ),
    .B2(_10324_),
    .C1(_10627_),
    .X(_10628_));
 sky130_fd_sc_hd__nor2_1 _14904_ (.A(_10069_),
    .B(_09760_),
    .Y(_10629_));
 sky130_fd_sc_hd__a22o_1 _14905_ (.A1(_10330_),
    .A2(\line_cache[129][1] ),
    .B1(\line_cache[128][1] ),
    .B2(_10629_),
    .X(_10630_));
 sky130_fd_sc_hd__a221o_1 _14906_ (.A1(\line_cache[131][1] ),
    .A2(_10328_),
    .B1(\line_cache[130][1] ),
    .B2(_10329_),
    .C1(_10630_),
    .X(_10631_));
 sky130_fd_sc_hd__a22o_1 _14907_ (.A1(_10336_),
    .A2(\line_cache[140][1] ),
    .B1(\line_cache[141][1] ),
    .B2(_10337_),
    .X(_10632_));
 sky130_fd_sc_hd__a221o_1 _14908_ (.A1(\line_cache[143][1] ),
    .A2(_10334_),
    .B1(\line_cache[142][1] ),
    .B2(_10335_),
    .C1(_10632_),
    .X(_10633_));
 sky130_fd_sc_hd__a22o_1 _14909_ (.A1(_10342_),
    .A2(\line_cache[139][1] ),
    .B1(\line_cache[138][1] ),
    .B2(_10343_),
    .X(_10634_));
 sky130_fd_sc_hd__a221o_1 _14910_ (.A1(\line_cache[137][1] ),
    .A2(_10340_),
    .B1(\line_cache[136][1] ),
    .B2(_10341_),
    .C1(_10634_),
    .X(_10635_));
 sky130_fd_sc_hd__or4_2 _14911_ (.A(_10628_),
    .B(_10631_),
    .C(_10633_),
    .D(_10635_),
    .X(_10636_));
 sky130_fd_sc_hd__nor2_1 _14912_ (.A(_10625_),
    .B(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__a22o_1 _14913_ (.A1(_10378_),
    .A2(\line_cache[80][1] ),
    .B1(_10379_),
    .B2(\line_cache[81][1] ),
    .X(_10638_));
 sky130_fd_sc_hd__a221o_1 _14914_ (.A1(\line_cache[83][1] ),
    .A2(_10376_),
    .B1(\line_cache[82][1] ),
    .B2(_10377_),
    .C1(_10638_),
    .X(_10639_));
 sky130_fd_sc_hd__a22o_1 _14915_ (.A1(_10384_),
    .A2(\line_cache[92][1] ),
    .B1(_10385_),
    .B2(\line_cache[93][1] ),
    .X(_10640_));
 sky130_fd_sc_hd__a221o_1 _14916_ (.A1(\line_cache[95][1] ),
    .A2(net136),
    .B1(\line_cache[94][1] ),
    .B2(_10383_),
    .C1(_10640_),
    .X(_10641_));
 sky130_fd_sc_hd__a22o_1 _14917_ (.A1(_10390_),
    .A2(\line_cache[84][1] ),
    .B1(_10391_),
    .B2(\line_cache[85][1] ),
    .X(_10642_));
 sky130_fd_sc_hd__a221o_1 _14918_ (.A1(\line_cache[87][1] ),
    .A2(_10388_),
    .B1(\line_cache[86][1] ),
    .B2(_10389_),
    .C1(_10642_),
    .X(_10643_));
 sky130_fd_sc_hd__a22o_1 _14919_ (.A1(_10396_),
    .A2(\line_cache[88][1] ),
    .B1(_10397_),
    .B2(\line_cache[89][1] ),
    .X(_10644_));
 sky130_fd_sc_hd__a221o_1 _14920_ (.A1(\line_cache[91][1] ),
    .A2(_10394_),
    .B1(\line_cache[90][1] ),
    .B2(_10395_),
    .C1(_10644_),
    .X(_10645_));
 sky130_fd_sc_hd__or4_1 _14921_ (.A(_10639_),
    .B(_10641_),
    .C(_10643_),
    .D(_10645_),
    .X(_10646_));
 sky130_fd_sc_hd__a22o_1 _14922_ (.A1(_10371_),
    .A2(\line_cache[100][1] ),
    .B1(_10372_),
    .B2(\line_cache[101][1] ),
    .X(_10647_));
 sky130_fd_sc_hd__a22o_1 _14923_ (.A1(_10369_),
    .A2(\line_cache[103][1] ),
    .B1(_10370_),
    .B2(\line_cache[102][1] ),
    .X(_10648_));
 sky130_fd_sc_hd__a22o_1 _14924_ (.A1(_10351_),
    .A2(\line_cache[96][1] ),
    .B1(_10352_),
    .B2(\line_cache[97][1] ),
    .X(_10649_));
 sky130_fd_sc_hd__a221o_1 _14925_ (.A1(\line_cache[99][1] ),
    .A2(_10349_),
    .B1(\line_cache[98][1] ),
    .B2(_10348_),
    .C1(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__clkbuf_4 _14926_ (.A(_10355_),
    .X(_10651_));
 sky130_fd_sc_hd__and3_1 _14927_ (.A(_10035_),
    .B(\line_cache[107][1] ),
    .C(_10651_),
    .X(_10652_));
 sky130_fd_sc_hd__and3_1 _14928_ (.A(_10176_),
    .B(\line_cache[105][1] ),
    .C(_10651_),
    .X(_10653_));
 sky130_fd_sc_hd__and3_1 _14929_ (.A(_10054_),
    .B(\line_cache[106][1] ),
    .C(_10651_),
    .X(_10654_));
 sky130_fd_sc_hd__and3_1 _14930_ (.A(_10360_),
    .B(\line_cache[104][1] ),
    .C(_10356_),
    .X(_10655_));
 sky130_fd_sc_hd__or4_1 _14931_ (.A(_10652_),
    .B(_10653_),
    .C(_10654_),
    .D(_10655_),
    .X(_10656_));
 sky130_fd_sc_hd__a22o_1 _14932_ (.A1(_10365_),
    .A2(\line_cache[108][1] ),
    .B1(_10366_),
    .B2(\line_cache[109][1] ),
    .X(_10657_));
 sky130_fd_sc_hd__a221o_1 _14933_ (.A1(\line_cache[111][1] ),
    .A2(_10363_),
    .B1(\line_cache[110][1] ),
    .B2(_10364_),
    .C1(_10657_),
    .X(_10658_));
 sky130_fd_sc_hd__or2_1 _14934_ (.A(_10656_),
    .B(_10658_),
    .X(_10659_));
 sky130_fd_sc_hd__or4_1 _14935_ (.A(_10647_),
    .B(_10648_),
    .C(_10650_),
    .D(_10659_),
    .X(_10660_));
 sky130_fd_sc_hd__nor2_1 _14936_ (.A(_10646_),
    .B(_10660_),
    .Y(_10661_));
 sky130_fd_sc_hd__and3_2 _14937_ (.A(_10613_),
    .B(_10637_),
    .C(_10661_),
    .X(_10662_));
 sky130_fd_sc_hd__nand3_1 _14938_ (.A(_10516_),
    .B(_10579_),
    .C(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__o21ba_2 _14939_ (.A1(_10405_),
    .A2(_10663_),
    .B1_N(_08979_),
    .X(_10664_));
 sky130_fd_sc_hd__buf_6 _14940_ (.A(_10664_),
    .X(net127));
 sky130_fd_sc_hd__and2b_1 _14941_ (.A_N(_09987_),
    .B(\line_cache[256][2] ),
    .X(_10665_));
 sky130_fd_sc_hd__and2b_1 _14942_ (.A_N(_09747_),
    .B(\line_cache[302][2] ),
    .X(_10666_));
 sky130_fd_sc_hd__a22o_1 _14943_ (.A1(_09743_),
    .A2(\line_cache[301][2] ),
    .B1(\line_cache[300][2] ),
    .B2(_09742_),
    .X(_10667_));
 sky130_fd_sc_hd__or3_1 _14944_ (.A(_10665_),
    .B(_10666_),
    .C(_10667_),
    .X(_10668_));
 sky130_fd_sc_hd__and3_1 _14945_ (.A(_09917_),
    .B(_09583_),
    .C(\line_cache[258][2] ),
    .X(_10669_));
 sky130_fd_sc_hd__and3_1 _14946_ (.A(_09848_),
    .B(_09583_),
    .C(\line_cache[260][2] ),
    .X(_10670_));
 sky130_fd_sc_hd__and3_1 _14947_ (.A(_09919_),
    .B(_09546_),
    .C(\line_cache[257][2] ),
    .X(_10671_));
 sky130_fd_sc_hd__and3_1 _14948_ (.A(_09840_),
    .B(_09546_),
    .C(\line_cache[259][2] ),
    .X(_10672_));
 sky130_fd_sc_hd__or4_1 _14949_ (.A(_10669_),
    .B(_10670_),
    .C(_10671_),
    .D(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__and3_1 _14950_ (.A(_09858_),
    .B(_09611_),
    .C(\line_cache[267][2] ),
    .X(_10674_));
 sky130_fd_sc_hd__a22o_1 _14951_ (.A1(_09998_),
    .A2(\line_cache[265][2] ),
    .B1(\line_cache[266][2] ),
    .B2(_09999_),
    .X(_10675_));
 sky130_fd_sc_hd__a311o_1 _14952_ (.A1(_09547_),
    .A2(\line_cache[268][2] ),
    .A3(_09862_),
    .B1(_10674_),
    .C1(_10675_),
    .X(_10676_));
 sky130_fd_sc_hd__nand2_1 _14953_ (.A(_10007_),
    .B(\line_cache[262][2] ),
    .Y(_10677_));
 sky130_fd_sc_hd__nand2_1 _14954_ (.A(_10010_),
    .B(\line_cache[261][2] ),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_1 _14955_ (.A(_10677_),
    .B(_10678_),
    .Y(_10679_));
 sky130_fd_sc_hd__a221oi_1 _14956_ (.A1(_10003_),
    .A2(\line_cache[264][2] ),
    .B1(_10005_),
    .B2(\line_cache[263][2] ),
    .C1(_10679_),
    .Y(_10680_));
 sky130_fd_sc_hd__or4b_1 _14957_ (.A(_10668_),
    .B(_10673_),
    .C(_10676_),
    .D_N(_10680_),
    .X(_10681_));
 sky130_fd_sc_hd__a22o_1 _14958_ (.A1(_09682_),
    .A2(\line_cache[308][2] ),
    .B1(\line_cache[309][2] ),
    .B2(_09685_),
    .X(_10682_));
 sky130_fd_sc_hd__a221o_1 _14959_ (.A1(\line_cache[311][2] ),
    .A2(_09689_),
    .B1(\line_cache[310][2] ),
    .B2(_09693_),
    .C1(_10682_),
    .X(_10683_));
 sky130_fd_sc_hd__a22o_1 _14960_ (.A1(_09728_),
    .A2(\line_cache[295][2] ),
    .B1(\line_cache[294][2] ),
    .B2(_09726_),
    .X(_10684_));
 sky130_fd_sc_hd__a221o_1 _14961_ (.A1(\line_cache[293][2] ),
    .A2(_09730_),
    .B1(\line_cache[292][2] ),
    .B2(_10018_),
    .C1(_10684_),
    .X(_10685_));
 sky130_fd_sc_hd__a22o_1 _14962_ (.A1(_09716_),
    .A2(\line_cache[296][2] ),
    .B1(\line_cache[297][2] ),
    .B2(_09721_),
    .X(_10686_));
 sky130_fd_sc_hd__a221o_1 _14963_ (.A1(\line_cache[299][2] ),
    .A2(_09718_),
    .B1(\line_cache[298][2] ),
    .B2(_09720_),
    .C1(_10686_),
    .X(_10687_));
 sky130_fd_sc_hd__a22o_1 _14964_ (.A1(_10025_),
    .A2(\line_cache[288][2] ),
    .B1(\line_cache[289][2] ),
    .B2(_10026_),
    .X(_10688_));
 sky130_fd_sc_hd__a221o_1 _14965_ (.A1(\line_cache[291][2] ),
    .A2(_10023_),
    .B1(\line_cache[290][2] ),
    .B2(_10024_),
    .C1(_10688_),
    .X(_10689_));
 sky130_fd_sc_hd__or4_2 _14966_ (.A(_10683_),
    .B(_10685_),
    .C(_10687_),
    .D(_10689_),
    .X(_10690_));
 sky130_fd_sc_hd__nor2_1 _14967_ (.A(_10681_),
    .B(_10690_),
    .Y(_10691_));
 sky130_fd_sc_hd__and3_1 _14968_ (.A(_10035_),
    .B(\line_cache[203][2] ),
    .C(_09538_),
    .X(_10692_));
 sky130_fd_sc_hd__and3_1 _14969_ (.A(_10038_),
    .B(\line_cache[206][2] ),
    .C(_09538_),
    .X(_10693_));
 sky130_fd_sc_hd__and3_1 _14970_ (.A(_10041_),
    .B(\line_cache[204][2] ),
    .C(_09539_),
    .X(_10694_));
 sky130_fd_sc_hd__a2111o_1 _14971_ (.A1(\line_cache[205][2] ),
    .A2(_10033_),
    .B1(_10692_),
    .C1(_10693_),
    .D1(_10694_),
    .X(_10695_));
 sky130_fd_sc_hd__a22o_1 _14972_ (.A1(_10049_),
    .A2(\line_cache[195][2] ),
    .B1(\line_cache[196][2] ),
    .B2(_10051_),
    .X(_10696_));
 sky130_fd_sc_hd__a221o_1 _14973_ (.A1(\line_cache[198][2] ),
    .A2(_10046_),
    .B1(\line_cache[197][2] ),
    .B2(_10047_),
    .C1(_10696_),
    .X(_10697_));
 sky130_fd_sc_hd__a22o_1 _14974_ (.A1(_10060_),
    .A2(\line_cache[200][2] ),
    .B1(_10063_),
    .B2(\line_cache[199][2] ),
    .X(_10698_));
 sky130_fd_sc_hd__a221o_1 _14975_ (.A1(\line_cache[202][2] ),
    .A2(_10056_),
    .B1(\line_cache[201][2] ),
    .B2(_10059_),
    .C1(_10698_),
    .X(_10699_));
 sky130_fd_sc_hd__and3_1 _14976_ (.A(_10067_),
    .B(\line_cache[193][2] ),
    .C(_09539_),
    .X(_10700_));
 sky130_fd_sc_hd__and3_1 _14977_ (.A(_10071_),
    .B(\line_cache[192][2] ),
    .C(_09539_),
    .X(_10701_));
 sky130_fd_sc_hd__and3_1 _14978_ (.A(_10074_),
    .B(\line_cache[194][2] ),
    .C(_09539_),
    .X(_10702_));
 sky130_fd_sc_hd__a2111o_1 _14979_ (.A1(_10066_),
    .A2(\line_cache[286][2] ),
    .B1(_10700_),
    .C1(_10701_),
    .D1(_10702_),
    .X(_10703_));
 sky130_fd_sc_hd__or4_1 _14980_ (.A(_10695_),
    .B(_10697_),
    .C(_10699_),
    .D(_10703_),
    .X(_10704_));
 sky130_fd_sc_hd__a22o_1 _14981_ (.A1(_09623_),
    .A2(\line_cache[275][2] ),
    .B1(_09620_),
    .B2(\line_cache[274][2] ),
    .X(_10705_));
 sky130_fd_sc_hd__a22o_1 _14982_ (.A1(_10080_),
    .A2(\line_cache[276][2] ),
    .B1(\line_cache[277][2] ),
    .B2(_10081_),
    .X(_10706_));
 sky130_fd_sc_hd__a22o_1 _14983_ (.A1(_10086_),
    .A2(\line_cache[270][2] ),
    .B1(\line_cache[269][2] ),
    .B2(_10088_),
    .X(_10707_));
 sky130_fd_sc_hd__a221o_1 _14984_ (.A1(\line_cache[273][2] ),
    .A2(_10083_),
    .B1(\line_cache[272][2] ),
    .B2(_10084_),
    .C1(_10707_),
    .X(_10708_));
 sky130_fd_sc_hd__a22o_1 _14985_ (.A1(_09655_),
    .A2(\line_cache[280][2] ),
    .B1(\line_cache[281][2] ),
    .B2(_09663_),
    .X(_10709_));
 sky130_fd_sc_hd__a22oi_1 _14986_ (.A1(_09661_),
    .A2(\line_cache[282][2] ),
    .B1(\line_cache[283][2] ),
    .B2(_09658_),
    .Y(_10710_));
 sky130_fd_sc_hd__a22oi_1 _14987_ (.A1(_09645_),
    .A2(\line_cache[285][2] ),
    .B1(\line_cache[284][2] ),
    .B2(_09648_),
    .Y(_10711_));
 sky130_fd_sc_hd__a22oi_1 _14988_ (.A1(_09636_),
    .A2(\line_cache[278][2] ),
    .B1(\line_cache[279][2] ),
    .B2(_09639_),
    .Y(_10712_));
 sky130_fd_sc_hd__and4b_1 _14989_ (.A_N(_10709_),
    .B(_10710_),
    .C(_10711_),
    .D(_10712_),
    .X(_10713_));
 sky130_fd_sc_hd__or4b_2 _14990_ (.A(_10705_),
    .B(_10706_),
    .C(_10708_),
    .D_N(_10713_),
    .X(_10714_));
 sky130_fd_sc_hd__nor2_1 _14991_ (.A(_10704_),
    .B(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__and3_1 _14992_ (.A(_10098_),
    .B(\line_cache[229][2] ),
    .C(_10100_),
    .X(_10716_));
 sky130_fd_sc_hd__and3_1 _14993_ (.A(_10102_),
    .B(\line_cache[230][2] ),
    .C(_10100_),
    .X(_10717_));
 sky130_fd_sc_hd__and3_1 _14994_ (.A(_10104_),
    .B(\line_cache[227][2] ),
    .C(_10100_),
    .X(_10718_));
 sky130_fd_sc_hd__and3_1 _14995_ (.A(_10106_),
    .B(\line_cache[228][2] ),
    .C(_10100_),
    .X(_10719_));
 sky130_fd_sc_hd__or4_1 _14996_ (.A(_10716_),
    .B(_10717_),
    .C(_10718_),
    .D(_10719_),
    .X(_10720_));
 sky130_fd_sc_hd__and3_1 _14997_ (.A(_09544_),
    .B(\line_cache[223][2] ),
    .C(_10109_),
    .X(_10721_));
 sky130_fd_sc_hd__and3_1 _14998_ (.A(_10071_),
    .B(\line_cache[224][2] ),
    .C(_10100_),
    .X(_10722_));
 sky130_fd_sc_hd__and3_1 _14999_ (.A(_10067_),
    .B(\line_cache[225][2] ),
    .C(_10100_),
    .X(_10723_));
 sky130_fd_sc_hd__and3_1 _15000_ (.A(_10074_),
    .B(\line_cache[226][2] ),
    .C(_10100_),
    .X(_10724_));
 sky130_fd_sc_hd__or4_1 _15001_ (.A(_10721_),
    .B(_10722_),
    .C(_10723_),
    .D(_10724_),
    .X(_10725_));
 sky130_fd_sc_hd__a22o_1 _15002_ (.A1(_10118_),
    .A2(\line_cache[236][2] ),
    .B1(_10120_),
    .B2(\line_cache[235][2] ),
    .X(_10726_));
 sky130_fd_sc_hd__a221o_1 _15003_ (.A1(\line_cache[238][2] ),
    .A2(_10116_),
    .B1(\line_cache[237][2] ),
    .B2(_10117_),
    .C1(_10726_),
    .X(_10727_));
 sky130_fd_sc_hd__a22o_1 _15004_ (.A1(_10125_),
    .A2(\line_cache[232][2] ),
    .B1(_10126_),
    .B2(\line_cache[231][2] ),
    .X(_10728_));
 sky130_fd_sc_hd__a221o_1 _15005_ (.A1(\line_cache[234][2] ),
    .A2(_10123_),
    .B1(\line_cache[233][2] ),
    .B2(_10124_),
    .C1(_10728_),
    .X(_10729_));
 sky130_fd_sc_hd__or4_1 _15006_ (.A(_10720_),
    .B(_10725_),
    .C(_10727_),
    .D(_10729_),
    .X(_10730_));
 sky130_fd_sc_hd__a22o_1 _15007_ (.A1(_10132_),
    .A2(\line_cache[220][2] ),
    .B1(_10133_),
    .B2(\line_cache[219][2] ),
    .X(_10731_));
 sky130_fd_sc_hd__a221o_1 _15008_ (.A1(\line_cache[222][2] ),
    .A2(_10130_),
    .B1(\line_cache[221][2] ),
    .B2(_10131_),
    .C1(_10731_),
    .X(_10732_));
 sky130_fd_sc_hd__a22o_1 _15009_ (.A1(_10138_),
    .A2(\line_cache[208][2] ),
    .B1(_10139_),
    .B2(\line_cache[207][2] ),
    .X(_10733_));
 sky130_fd_sc_hd__a221o_1 _15010_ (.A1(\line_cache[210][2] ),
    .A2(_10136_),
    .B1(\line_cache[209][2] ),
    .B2(_10137_),
    .C1(_10733_),
    .X(_10734_));
 sky130_fd_sc_hd__a22o_1 _15011_ (.A1(_10144_),
    .A2(\line_cache[216][2] ),
    .B1(_10145_),
    .B2(\line_cache[215][2] ),
    .X(_10735_));
 sky130_fd_sc_hd__a221o_1 _15012_ (.A1(\line_cache[218][2] ),
    .A2(_10142_),
    .B1(\line_cache[217][2] ),
    .B2(_10143_),
    .C1(_10735_),
    .X(_10736_));
 sky130_fd_sc_hd__and2b_1 _15013_ (.A_N(_10148_),
    .B(\line_cache[211][2] ),
    .X(_10737_));
 sky130_fd_sc_hd__and2b_1 _15014_ (.A_N(_10150_),
    .B(\line_cache[212][2] ),
    .X(_10738_));
 sky130_fd_sc_hd__and2b_1 _15015_ (.A_N(_10152_),
    .B(\line_cache[213][2] ),
    .X(_10739_));
 sky130_fd_sc_hd__and2b_1 _15016_ (.A_N(_10154_),
    .B(\line_cache[214][2] ),
    .X(_10740_));
 sky130_fd_sc_hd__or4_1 _15017_ (.A(_10737_),
    .B(_10738_),
    .C(_10739_),
    .D(_10740_),
    .X(_10741_));
 sky130_fd_sc_hd__or4_2 _15018_ (.A(_10732_),
    .B(_10734_),
    .C(_10736_),
    .D(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(_10730_),
    .B(_10742_),
    .Y(_10743_));
 sky130_fd_sc_hd__and3_1 _15020_ (.A(_10031_),
    .B(\line_cache[77][2] ),
    .C(_10167_),
    .X(_10744_));
 sky130_fd_sc_hd__and3_1 _15021_ (.A(_10038_),
    .B(\line_cache[78][2] ),
    .C(_10161_),
    .X(_10745_));
 sky130_fd_sc_hd__and3_1 _15022_ (.A(_10041_),
    .B(\line_cache[76][2] ),
    .C(_10161_),
    .X(_10746_));
 sky130_fd_sc_hd__a2111o_1 _15023_ (.A1(_10168_),
    .A2(\line_cache[79][2] ),
    .B1(_10744_),
    .C1(_10745_),
    .D1(_10746_),
    .X(_10747_));
 sky130_fd_sc_hd__a22o_1 _15024_ (.A1(_10182_),
    .A2(\line_cache[64][2] ),
    .B1(_10183_),
    .B2(\line_cache[65][2] ),
    .X(_10748_));
 sky130_fd_sc_hd__a221o_1 _15025_ (.A1(\line_cache[67][2] ),
    .A2(_10180_),
    .B1(\line_cache[66][2] ),
    .B2(_10181_),
    .C1(_10748_),
    .X(_10749_));
 sky130_fd_sc_hd__nor2_2 _15026_ (.A(_09766_),
    .B(_10045_),
    .Y(_10750_));
 sky130_fd_sc_hd__a22o_1 _15027_ (.A1(_10163_),
    .A2(\line_cache[68][2] ),
    .B1(_10164_),
    .B2(\line_cache[69][2] ),
    .X(_10751_));
 sky130_fd_sc_hd__a221o_1 _15028_ (.A1(\line_cache[71][2] ),
    .A2(_10159_),
    .B1(\line_cache[70][2] ),
    .B2(_10750_),
    .C1(_10751_),
    .X(_10752_));
 sky130_fd_sc_hd__nor2_1 _15029_ (.A(_09766_),
    .B(_10058_),
    .Y(_10753_));
 sky130_fd_sc_hd__a22o_1 _15030_ (.A1(_10175_),
    .A2(\line_cache[72][2] ),
    .B1(_10753_),
    .B2(\line_cache[73][2] ),
    .X(_10754_));
 sky130_fd_sc_hd__a221o_1 _15031_ (.A1(\line_cache[75][2] ),
    .A2(_10173_),
    .B1(\line_cache[74][2] ),
    .B2(_10174_),
    .C1(_10754_),
    .X(_10755_));
 sky130_fd_sc_hd__or4_4 _15032_ (.A(_10747_),
    .B(_10749_),
    .C(_10752_),
    .D(_10755_),
    .X(_10756_));
 sky130_fd_sc_hd__a22o_1 _15033_ (.A1(_10189_),
    .A2(\line_cache[252][2] ),
    .B1(_10190_),
    .B2(\line_cache[251][2] ),
    .X(_10757_));
 sky130_fd_sc_hd__a221o_1 _15034_ (.A1(\line_cache[254][2] ),
    .A2(_10187_),
    .B1(\line_cache[253][2] ),
    .B2(_10188_),
    .C1(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__a22o_1 _15035_ (.A1(_10195_),
    .A2(\line_cache[248][2] ),
    .B1(_10196_),
    .B2(\line_cache[247][2] ),
    .X(_10759_));
 sky130_fd_sc_hd__a221o_1 _15036_ (.A1(\line_cache[250][2] ),
    .A2(_10193_),
    .B1(\line_cache[249][2] ),
    .B2(_10194_),
    .C1(_10759_),
    .X(_10760_));
 sky130_fd_sc_hd__and2b_1 _15037_ (.A_N(_10200_),
    .B(\line_cache[240][2] ),
    .X(_10761_));
 sky130_fd_sc_hd__and2b_1 _15038_ (.A_N(_09570_),
    .B(\line_cache[241][2] ),
    .X(_10762_));
 sky130_fd_sc_hd__and2b_1 _15039_ (.A_N(_10203_),
    .B(\line_cache[242][2] ),
    .X(_10763_));
 sky130_fd_sc_hd__a2111o_1 _15040_ (.A1(\line_cache[239][2] ),
    .A2(_10199_),
    .B1(_10761_),
    .C1(_10762_),
    .D1(_10763_),
    .X(_10764_));
 sky130_fd_sc_hd__and2b_1 _15041_ (.A_N(_10206_),
    .B(\line_cache[243][2] ),
    .X(_10765_));
 sky130_fd_sc_hd__and2b_1 _15042_ (.A_N(_10208_),
    .B(\line_cache[244][2] ),
    .X(_10766_));
 sky130_fd_sc_hd__and2b_1 _15043_ (.A_N(_09597_),
    .B(\line_cache[245][2] ),
    .X(_10767_));
 sky130_fd_sc_hd__and2b_1 _15044_ (.A_N(_10211_),
    .B(\line_cache[246][2] ),
    .X(_10768_));
 sky130_fd_sc_hd__or4_1 _15045_ (.A(_10765_),
    .B(_10766_),
    .C(_10767_),
    .D(_10768_),
    .X(_10769_));
 sky130_fd_sc_hd__or4_1 _15046_ (.A(_10758_),
    .B(_10760_),
    .C(_10764_),
    .D(_10769_),
    .X(_10770_));
 sky130_fd_sc_hd__nor2_1 _15047_ (.A(_10756_),
    .B(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__and4_2 _15048_ (.A(_10691_),
    .B(_10715_),
    .C(_10743_),
    .D(_10771_),
    .X(_10772_));
 sky130_fd_sc_hd__a22o_1 _15049_ (.A1(_09842_),
    .A2(\line_cache[6][2] ),
    .B1(\line_cache[5][2] ),
    .B2(_09844_),
    .X(_10773_));
 sky130_fd_sc_hd__a221o_1 _15050_ (.A1(\line_cache[4][2] ),
    .A2(_09850_),
    .B1(\line_cache[3][2] ),
    .B2(_09914_),
    .C1(_10773_),
    .X(_10774_));
 sky130_fd_sc_hd__and3_1 _15051_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][2] ),
    .X(_10775_));
 sky130_fd_sc_hd__and3_1 _15052_ (.A(_09919_),
    .B(_09532_),
    .C(\line_cache[1][2] ),
    .X(_10776_));
 sky130_fd_sc_hd__a211o_1 _15053_ (.A1(\line_cache[15][2] ),
    .A2(_09867_),
    .B1(_10775_),
    .C1(_10776_),
    .X(_10777_));
 sky130_fd_sc_hd__and3_1 _15054_ (.A(_09922_),
    .B(_09531_),
    .C(\line_cache[63][2] ),
    .X(_10778_));
 sky130_fd_sc_hd__a31o_1 _15055_ (.A1(_09547_),
    .A2(\line_cache[319][2] ),
    .A3(_09922_),
    .B1(_10778_),
    .X(_10779_));
 sky130_fd_sc_hd__a221o_1 _15056_ (.A1(\line_cache[47][2] ),
    .A2(_09806_),
    .B1(\line_cache[31][2] ),
    .B2(_09907_),
    .C1(_10779_),
    .X(_10780_));
 sky130_fd_sc_hd__nand2_1 _15057_ (.A(_09746_),
    .B(\line_cache[303][2] ),
    .Y(_10781_));
 sky130_fd_sc_hd__nand2_1 _15058_ (.A(_09930_),
    .B(\line_cache[271][2] ),
    .Y(_10782_));
 sky130_fd_sc_hd__nand2_1 _15059_ (.A(_10781_),
    .B(_10782_),
    .Y(_10783_));
 sky130_fd_sc_hd__a221oi_2 _15060_ (.A1(\line_cache[255][2] ),
    .A2(_09926_),
    .B1(\line_cache[287][2] ),
    .B2(_09927_),
    .C1(_10783_),
    .Y(_10784_));
 sky130_fd_sc_hd__or4b_1 _15061_ (.A(_10774_),
    .B(_10777_),
    .C(_10780_),
    .D_N(_10784_),
    .X(_10785_));
 sky130_fd_sc_hd__a22o_1 _15062_ (.A1(_09803_),
    .A2(\line_cache[45][2] ),
    .B1(\line_cache[46][2] ),
    .B2(_09804_),
    .X(_10786_));
 sky130_fd_sc_hd__a22o_1 _15063_ (.A1(_09824_),
    .A2(\line_cache[48][2] ),
    .B1(\line_cache[49][2] ),
    .B2(_09826_),
    .X(_10787_));
 sky130_fd_sc_hd__nand2_1 _15064_ (.A(_09787_),
    .B(\line_cache[41][2] ),
    .Y(_10788_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(_09789_),
    .B(\line_cache[42][2] ),
    .Y(_10789_));
 sky130_fd_sc_hd__nand2_1 _15066_ (.A(_10788_),
    .B(_10789_),
    .Y(_10790_));
 sky130_fd_sc_hd__a221oi_4 _15067_ (.A1(_09785_),
    .A2(\line_cache[43][2] ),
    .B1(\line_cache[44][2] ),
    .B2(_09801_),
    .C1(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__or3b_1 _15068_ (.A(_10786_),
    .B(_10787_),
    .C_N(_10791_),
    .X(_10792_));
 sky130_fd_sc_hd__a22o_1 _15069_ (.A1(_09699_),
    .A2(\line_cache[317][2] ),
    .B1(\line_cache[316][2] ),
    .B2(_09697_),
    .X(_10793_));
 sky130_fd_sc_hd__a22o_1 _15070_ (.A1(_09832_),
    .A2(\line_cache[58][2] ),
    .B1(\line_cache[59][2] ),
    .B2(_09833_),
    .X(_10794_));
 sky130_fd_sc_hd__a22o_1 _15071_ (.A1(_09819_),
    .A2(\line_cache[61][2] ),
    .B1(\line_cache[60][2] ),
    .B2(_09817_),
    .X(_10795_));
 sky130_fd_sc_hd__a22o_1 _15072_ (.A1(_09822_),
    .A2(\line_cache[62][2] ),
    .B1(\line_cache[318][2] ),
    .B2(_09702_),
    .X(_10796_));
 sky130_fd_sc_hd__or4_1 _15073_ (.A(_10793_),
    .B(_10794_),
    .C(_10795_),
    .D(_10796_),
    .X(_10797_));
 sky130_fd_sc_hd__a22o_1 _15074_ (.A1(_09675_),
    .A2(\line_cache[304][2] ),
    .B1(\line_cache[305][2] ),
    .B2(_09676_),
    .X(_10798_));
 sky130_fd_sc_hd__a22o_1 _15075_ (.A1(_09705_),
    .A2(\line_cache[312][2] ),
    .B1(\line_cache[313][2] ),
    .B2(_09707_),
    .X(_10799_));
 sky130_fd_sc_hd__a22o_1 _15076_ (.A1(_09708_),
    .A2(\line_cache[314][2] ),
    .B1(\line_cache[315][2] ),
    .B2(_09709_),
    .X(_10800_));
 sky130_fd_sc_hd__a22o_1 _15077_ (.A1(_09677_),
    .A2(\line_cache[306][2] ),
    .B1(\line_cache[307][2] ),
    .B2(_09678_),
    .X(_10801_));
 sky130_fd_sc_hd__or4_1 _15078_ (.A(_10798_),
    .B(_10799_),
    .C(_10800_),
    .D(_10801_),
    .X(_10802_));
 sky130_fd_sc_hd__a22o_1 _15079_ (.A1(_09830_),
    .A2(\line_cache[56][2] ),
    .B1(\line_cache[57][2] ),
    .B2(_09834_),
    .X(_10803_));
 sky130_fd_sc_hd__a22o_1 _15080_ (.A1(_09809_),
    .A2(\line_cache[52][2] ),
    .B1(\line_cache[53][2] ),
    .B2(_09811_),
    .X(_10804_));
 sky130_fd_sc_hd__a22o_1 _15081_ (.A1(_09827_),
    .A2(\line_cache[50][2] ),
    .B1(\line_cache[51][2] ),
    .B2(_09828_),
    .X(_10805_));
 sky130_fd_sc_hd__a22o_1 _15082_ (.A1(_09813_),
    .A2(\line_cache[54][2] ),
    .B1(\line_cache[55][2] ),
    .B2(_09815_),
    .X(_10806_));
 sky130_fd_sc_hd__or4_1 _15083_ (.A(_10803_),
    .B(_10804_),
    .C(_10805_),
    .D(_10806_),
    .X(_10807_));
 sky130_fd_sc_hd__or4_2 _15084_ (.A(_10792_),
    .B(_10797_),
    .C(_10802_),
    .D(_10807_),
    .X(_10808_));
 sky130_fd_sc_hd__nand2_1 _15085_ (.A(_09864_),
    .B(\line_cache[12][2] ),
    .Y(_10809_));
 sky130_fd_sc_hd__nand2_1 _15086_ (.A(_09860_),
    .B(\line_cache[11][2] ),
    .Y(_10810_));
 sky130_fd_sc_hd__nand2_1 _15087_ (.A(_10809_),
    .B(_10810_),
    .Y(_10811_));
 sky130_fd_sc_hd__a221oi_2 _15088_ (.A1(_09870_),
    .A2(\line_cache[14][2] ),
    .B1(\line_cache[13][2] ),
    .B2(_09873_),
    .C1(_10811_),
    .Y(_10812_));
 sky130_fd_sc_hd__nand2_1 _15089_ (.A(_09853_),
    .B(\line_cache[10][2] ),
    .Y(_10813_));
 sky130_fd_sc_hd__nand2_1 _15090_ (.A(_09857_),
    .B(\line_cache[9][2] ),
    .Y(_10814_));
 sky130_fd_sc_hd__nand2_1 _15091_ (.A(_10813_),
    .B(_10814_),
    .Y(_10815_));
 sky130_fd_sc_hd__a221oi_1 _15092_ (.A1(_09855_),
    .A2(\line_cache[8][2] ),
    .B1(_09847_),
    .B2(\line_cache[7][2] ),
    .C1(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__nand2_1 _15093_ (.A(_10812_),
    .B(_10816_),
    .Y(_10817_));
 sky130_fd_sc_hd__and3_1 _15094_ (.A(_09631_),
    .B(_09532_),
    .C(\line_cache[21][2] ),
    .X(_10818_));
 sky130_fd_sc_hd__a22o_1 _15095_ (.A1(_09884_),
    .A2(\line_cache[23][2] ),
    .B1(\line_cache[22][2] ),
    .B2(_09886_),
    .X(_10819_));
 sky130_fd_sc_hd__a22o_1 _15096_ (.A1(_09877_),
    .A2(\line_cache[19][2] ),
    .B1(\line_cache[18][2] ),
    .B2(_09878_),
    .X(_10820_));
 sky130_fd_sc_hd__a221o_1 _15097_ (.A1(\line_cache[17][2] ),
    .A2(_09969_),
    .B1(\line_cache[16][2] ),
    .B2(_09970_),
    .C1(_10820_),
    .X(_10821_));
 sky130_fd_sc_hd__a2111o_1 _15098_ (.A1(\line_cache[20][2] ),
    .A2(_09888_),
    .B1(_10818_),
    .C1(_10819_),
    .D1(_10821_),
    .X(_10822_));
 sky130_fd_sc_hd__a22o_1 _15099_ (.A1(_09890_),
    .A2(\line_cache[27][2] ),
    .B1(\line_cache[26][2] ),
    .B2(_09896_),
    .X(_10823_));
 sky130_fd_sc_hd__a221o_1 _15100_ (.A1(\line_cache[25][2] ),
    .A2(_09892_),
    .B1(\line_cache[24][2] ),
    .B2(_09895_),
    .C1(_10823_),
    .X(_10824_));
 sky130_fd_sc_hd__a22o_1 _15101_ (.A1(_09796_),
    .A2(\line_cache[33][2] ),
    .B1(\line_cache[34][2] ),
    .B2(_09798_),
    .X(_10825_));
 sky130_fd_sc_hd__a221oi_1 _15102_ (.A1(\line_cache[36][2] ),
    .A2(_09777_),
    .B1(\line_cache[35][2] ),
    .B2(_09794_),
    .C1(_10825_),
    .Y(_10826_));
 sky130_fd_sc_hd__nand2_1 _15103_ (.A(_09773_),
    .B(\line_cache[38][2] ),
    .Y(_10827_));
 sky130_fd_sc_hd__nand2_1 _15104_ (.A(_09775_),
    .B(\line_cache[37][2] ),
    .Y(_10828_));
 sky130_fd_sc_hd__nand2_1 _15105_ (.A(_10827_),
    .B(_10828_),
    .Y(_10829_));
 sky130_fd_sc_hd__a221oi_1 _15106_ (.A1(_09783_),
    .A2(\line_cache[40][2] ),
    .B1(\line_cache[39][2] ),
    .B2(_09780_),
    .C1(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__nand2_1 _15107_ (.A(_10826_),
    .B(_10830_),
    .Y(_10831_));
 sky130_fd_sc_hd__a22o_1 _15108_ (.A1(_09903_),
    .A2(\line_cache[29][2] ),
    .B1(\line_cache[28][2] ),
    .B2(_09900_),
    .X(_10832_));
 sky130_fd_sc_hd__a221o_1 _15109_ (.A1(\line_cache[32][2] ),
    .A2(_09792_),
    .B1(\line_cache[30][2] ),
    .B2(_09905_),
    .C1(_10832_),
    .X(_10833_));
 sky130_fd_sc_hd__nor3_1 _15110_ (.A(_10824_),
    .B(_10831_),
    .C(_10833_),
    .Y(_10834_));
 sky130_fd_sc_hd__or3b_1 _15111_ (.A(_10817_),
    .B(_10822_),
    .C_N(_10834_),
    .X(_10835_));
 sky130_fd_sc_hd__nor3_1 _15112_ (.A(_10785_),
    .B(_10808_),
    .C(_10835_),
    .Y(_10836_));
 sky130_fd_sc_hd__a22o_1 _15113_ (.A1(_10390_),
    .A2(\line_cache[84][2] ),
    .B1(_10391_),
    .B2(\line_cache[85][2] ),
    .X(_10837_));
 sky130_fd_sc_hd__a22o_1 _15114_ (.A1(_10388_),
    .A2(\line_cache[87][2] ),
    .B1(_10389_),
    .B2(\line_cache[86][2] ),
    .X(_10838_));
 sky130_fd_sc_hd__or2_1 _15115_ (.A(_10837_),
    .B(_10838_),
    .X(_10839_));
 sky130_fd_sc_hd__a22o_1 _15116_ (.A1(_10378_),
    .A2(\line_cache[80][2] ),
    .B1(_10379_),
    .B2(\line_cache[81][2] ),
    .X(_10840_));
 sky130_fd_sc_hd__a221o_1 _15117_ (.A1(\line_cache[83][2] ),
    .A2(_10376_),
    .B1(\line_cache[82][2] ),
    .B2(_10377_),
    .C1(_10840_),
    .X(_10841_));
 sky130_fd_sc_hd__a22o_1 _15118_ (.A1(_10384_),
    .A2(\line_cache[92][2] ),
    .B1(_10385_),
    .B2(\line_cache[93][2] ),
    .X(_10842_));
 sky130_fd_sc_hd__a221o_1 _15119_ (.A1(\line_cache[95][2] ),
    .A2(net136),
    .B1(\line_cache[94][2] ),
    .B2(_10383_),
    .C1(_10842_),
    .X(_10843_));
 sky130_fd_sc_hd__a22o_1 _15120_ (.A1(_10396_),
    .A2(\line_cache[88][2] ),
    .B1(_10397_),
    .B2(\line_cache[89][2] ),
    .X(_10844_));
 sky130_fd_sc_hd__a221o_1 _15121_ (.A1(\line_cache[91][2] ),
    .A2(_10394_),
    .B1(\line_cache[90][2] ),
    .B2(_10395_),
    .C1(_10844_),
    .X(_10845_));
 sky130_fd_sc_hd__or4_2 _15122_ (.A(_10839_),
    .B(_10841_),
    .C(_10843_),
    .D(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__a22o_1 _15123_ (.A1(_10371_),
    .A2(\line_cache[100][2] ),
    .B1(_10372_),
    .B2(\line_cache[101][2] ),
    .X(_10847_));
 sky130_fd_sc_hd__a22o_1 _15124_ (.A1(_10369_),
    .A2(\line_cache[103][2] ),
    .B1(_10370_),
    .B2(\line_cache[102][2] ),
    .X(_10848_));
 sky130_fd_sc_hd__a22o_1 _15125_ (.A1(_10351_),
    .A2(\line_cache[96][2] ),
    .B1(_10352_),
    .B2(\line_cache[97][2] ),
    .X(_10849_));
 sky130_fd_sc_hd__a221o_2 _15126_ (.A1(\line_cache[99][2] ),
    .A2(_10349_),
    .B1(\line_cache[98][2] ),
    .B2(_10348_),
    .C1(_10849_),
    .X(_10850_));
 sky130_fd_sc_hd__and3_1 _15127_ (.A(_10035_),
    .B(\line_cache[107][2] ),
    .C(_10355_),
    .X(_10851_));
 sky130_fd_sc_hd__and3_1 _15128_ (.A(_10176_),
    .B(\line_cache[105][2] ),
    .C(_10651_),
    .X(_10852_));
 sky130_fd_sc_hd__and3_1 _15129_ (.A(_10054_),
    .B(\line_cache[106][2] ),
    .C(_10651_),
    .X(_10853_));
 sky130_fd_sc_hd__and3_1 _15130_ (.A(_10360_),
    .B(\line_cache[104][2] ),
    .C(_10651_),
    .X(_10854_));
 sky130_fd_sc_hd__or4_1 _15131_ (.A(_10851_),
    .B(_10852_),
    .C(_10853_),
    .D(_10854_),
    .X(_10855_));
 sky130_fd_sc_hd__a22o_1 _15132_ (.A1(_10365_),
    .A2(\line_cache[108][2] ),
    .B1(_10366_),
    .B2(\line_cache[109][2] ),
    .X(_10856_));
 sky130_fd_sc_hd__a221o_1 _15133_ (.A1(\line_cache[111][2] ),
    .A2(_10363_),
    .B1(\line_cache[110][2] ),
    .B2(_10364_),
    .C1(_10856_),
    .X(_10857_));
 sky130_fd_sc_hd__or2_1 _15134_ (.A(_10855_),
    .B(_10857_),
    .X(_10858_));
 sky130_fd_sc_hd__or4_1 _15135_ (.A(_10847_),
    .B(_10848_),
    .C(_10850_),
    .D(_10858_),
    .X(_10859_));
 sky130_fd_sc_hd__nor2_1 _15136_ (.A(_10846_),
    .B(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__a22o_1 _15137_ (.A1(_10219_),
    .A2(\line_cache[157][2] ),
    .B1(\line_cache[156][2] ),
    .B2(_10220_),
    .X(_10861_));
 sky130_fd_sc_hd__a221o_1 _15138_ (.A1(\line_cache[159][2] ),
    .A2(_10217_),
    .B1(\line_cache[158][2] ),
    .B2(_10218_),
    .C1(_10861_),
    .X(_10862_));
 sky130_fd_sc_hd__a22o_1 _15139_ (.A1(_10231_),
    .A2(\line_cache[147][2] ),
    .B1(\line_cache[146][2] ),
    .B2(_10232_),
    .X(_10863_));
 sky130_fd_sc_hd__a221oi_2 _15140_ (.A1(\line_cache[145][2] ),
    .A2(_10229_),
    .B1(\line_cache[144][2] ),
    .B2(_10230_),
    .C1(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__a22o_1 _15141_ (.A1(_10225_),
    .A2(\line_cache[151][2] ),
    .B1(\line_cache[150][2] ),
    .B2(_10226_),
    .X(_10865_));
 sky130_fd_sc_hd__a221oi_2 _15142_ (.A1(\line_cache[149][2] ),
    .A2(_10223_),
    .B1(\line_cache[148][2] ),
    .B2(_10224_),
    .C1(_10865_),
    .Y(_10866_));
 sky130_fd_sc_hd__a22o_1 _15143_ (.A1(_10237_),
    .A2(\line_cache[155][2] ),
    .B1(\line_cache[154][2] ),
    .B2(_10238_),
    .X(_10867_));
 sky130_fd_sc_hd__a221oi_2 _15144_ (.A1(\line_cache[153][2] ),
    .A2(_10235_),
    .B1(\line_cache[152][2] ),
    .B2(_10236_),
    .C1(_10867_),
    .Y(_10868_));
 sky130_fd_sc_hd__and4b_1 _15145_ (.A_N(_10862_),
    .B(_10864_),
    .C(_10866_),
    .D(_10868_),
    .X(_10869_));
 sky130_fd_sc_hd__a22o_1 _15146_ (.A1(_10244_),
    .A2(\line_cache[173][2] ),
    .B1(\line_cache[172][2] ),
    .B2(_10245_),
    .X(_10870_));
 sky130_fd_sc_hd__a221o_1 _15147_ (.A1(\line_cache[175][2] ),
    .A2(_10242_),
    .B1(\line_cache[174][2] ),
    .B2(_10243_),
    .C1(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__a22o_1 _15148_ (.A1(_10250_),
    .A2(\line_cache[165][2] ),
    .B1(\line_cache[164][2] ),
    .B2(_10251_),
    .X(_10872_));
 sky130_fd_sc_hd__a221oi_1 _15149_ (.A1(\line_cache[167][2] ),
    .A2(_10248_),
    .B1(\line_cache[166][2] ),
    .B2(_10249_),
    .C1(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__a22o_1 _15150_ (.A1(_10256_),
    .A2(\line_cache[160][2] ),
    .B1(\line_cache[161][2] ),
    .B2(_10257_),
    .X(_10874_));
 sky130_fd_sc_hd__a221oi_2 _15151_ (.A1(\line_cache[163][2] ),
    .A2(_10254_),
    .B1(\line_cache[162][2] ),
    .B2(_10255_),
    .C1(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__a22o_1 _15152_ (.A1(_10261_),
    .A2(\line_cache[168][2] ),
    .B1(\line_cache[169][2] ),
    .B2(_10260_),
    .X(_10876_));
 sky130_fd_sc_hd__a221oi_4 _15153_ (.A1(\line_cache[171][2] ),
    .A2(_10262_),
    .B1(\line_cache[170][2] ),
    .B2(_10263_),
    .C1(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__and4b_1 _15154_ (.A_N(_10871_),
    .B(_10873_),
    .C(_10875_),
    .D(_10877_),
    .X(_10878_));
 sky130_fd_sc_hd__a22o_1 _15155_ (.A1(_10277_),
    .A2(\line_cache[184][2] ),
    .B1(\line_cache[185][2] ),
    .B2(_10278_),
    .X(_10879_));
 sky130_fd_sc_hd__a221o_1 _15156_ (.A1(\line_cache[187][2] ),
    .A2(_10275_),
    .B1(\line_cache[186][2] ),
    .B2(_10276_),
    .C1(_10879_),
    .X(_10880_));
 sky130_fd_sc_hd__a22o_1 _15157_ (.A1(_10284_),
    .A2(\line_cache[176][2] ),
    .B1(_10285_),
    .B2(\line_cache[177][2] ),
    .X(_10881_));
 sky130_fd_sc_hd__a221oi_2 _15158_ (.A1(\line_cache[179][2] ),
    .A2(_10282_),
    .B1(\line_cache[178][2] ),
    .B2(_10283_),
    .C1(_10881_),
    .Y(_10882_));
 sky130_fd_sc_hd__and3_1 _15159_ (.A(_10288_),
    .B(_10102_),
    .C(\line_cache[182][2] ),
    .X(_10883_));
 sky130_fd_sc_hd__and3_1 _15160_ (.A(_09755_),
    .B(_10098_),
    .C(\line_cache[181][2] ),
    .X(_10884_));
 sky130_fd_sc_hd__a31o_1 _15161_ (.A1(\line_cache[180][2] ),
    .A2(_10288_),
    .A3(_10106_),
    .B1(_10884_),
    .X(_10885_));
 sky130_fd_sc_hd__a311oi_2 _15162_ (.A1(\line_cache[183][2] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_10883_),
    .C1(_10885_),
    .Y(_10886_));
 sky130_fd_sc_hd__a22o_1 _15163_ (.A1(_10272_),
    .A2(\line_cache[189][2] ),
    .B1(\line_cache[188][2] ),
    .B2(_10271_),
    .X(_10887_));
 sky130_fd_sc_hd__a221oi_1 _15164_ (.A1(\line_cache[191][2] ),
    .A2(_10269_),
    .B1(\line_cache[190][2] ),
    .B2(_10270_),
    .C1(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__and4b_1 _15165_ (.A_N(_10880_),
    .B(_10882_),
    .C(_10886_),
    .D(_10888_),
    .X(_10889_));
 sky130_fd_sc_hd__and3_2 _15166_ (.A(_10869_),
    .B(_10878_),
    .C(_10889_),
    .X(_10890_));
 sky130_fd_sc_hd__a22o_1 _15167_ (.A1(_10298_),
    .A2(\line_cache[112][2] ),
    .B1(_10299_),
    .B2(\line_cache[113][2] ),
    .X(_10891_));
 sky130_fd_sc_hd__a221o_1 _15168_ (.A1(\line_cache[115][2] ),
    .A2(_10296_),
    .B1(\line_cache[114][2] ),
    .B2(_10297_),
    .C1(_10891_),
    .X(_10892_));
 sky130_fd_sc_hd__a22o_1 _15169_ (.A1(_10305_),
    .A2(\line_cache[124][2] ),
    .B1(_10306_),
    .B2(\line_cache[125][2] ),
    .X(_10893_));
 sky130_fd_sc_hd__a221o_1 _15170_ (.A1(\line_cache[127][2] ),
    .A2(_10303_),
    .B1(\line_cache[126][2] ),
    .B2(_10304_),
    .C1(_10893_),
    .X(_10894_));
 sky130_fd_sc_hd__a22o_1 _15171_ (.A1(_10311_),
    .A2(\line_cache[116][2] ),
    .B1(_10312_),
    .B2(\line_cache[117][2] ),
    .X(_10895_));
 sky130_fd_sc_hd__a221o_1 _15172_ (.A1(\line_cache[119][2] ),
    .A2(_10309_),
    .B1(\line_cache[118][2] ),
    .B2(_10310_),
    .C1(_10895_),
    .X(_10896_));
 sky130_fd_sc_hd__a22o_1 _15173_ (.A1(_10317_),
    .A2(\line_cache[120][2] ),
    .B1(_10318_),
    .B2(\line_cache[121][2] ),
    .X(_10897_));
 sky130_fd_sc_hd__a221o_1 _15174_ (.A1(\line_cache[123][2] ),
    .A2(_10315_),
    .B1(\line_cache[122][2] ),
    .B2(_10316_),
    .C1(_10897_),
    .X(_10898_));
 sky130_fd_sc_hd__or4_1 _15175_ (.A(_10892_),
    .B(_10894_),
    .C(_10896_),
    .D(_10898_),
    .X(_10899_));
 sky130_fd_sc_hd__and3_1 _15176_ (.A(_09758_),
    .B(_10098_),
    .C(\line_cache[133][2] ),
    .X(_10900_));
 sky130_fd_sc_hd__a21o_1 _15177_ (.A1(\line_cache[132][2] ),
    .A2(_10324_),
    .B1(_10900_),
    .X(_10901_));
 sky130_fd_sc_hd__a221o_1 _15178_ (.A1(\line_cache[135][2] ),
    .A2(_10322_),
    .B1(\line_cache[134][2] ),
    .B2(_10323_),
    .C1(_10901_),
    .X(_10902_));
 sky130_fd_sc_hd__and3_1 _15179_ (.A(_10071_),
    .B(\line_cache[128][2] ),
    .C(_09758_),
    .X(_10903_));
 sky130_fd_sc_hd__a21o_1 _15180_ (.A1(\line_cache[129][2] ),
    .A2(_10330_),
    .B1(_10903_),
    .X(_10904_));
 sky130_fd_sc_hd__a221o_1 _15181_ (.A1(\line_cache[131][2] ),
    .A2(_10328_),
    .B1(\line_cache[130][2] ),
    .B2(_10329_),
    .C1(_10904_),
    .X(_10905_));
 sky130_fd_sc_hd__a22o_1 _15182_ (.A1(_10336_),
    .A2(\line_cache[140][2] ),
    .B1(\line_cache[141][2] ),
    .B2(_10337_),
    .X(_10906_));
 sky130_fd_sc_hd__a221o_1 _15183_ (.A1(\line_cache[143][2] ),
    .A2(_10334_),
    .B1(\line_cache[142][2] ),
    .B2(_10335_),
    .C1(_10906_),
    .X(_10907_));
 sky130_fd_sc_hd__a22o_1 _15184_ (.A1(_10342_),
    .A2(\line_cache[139][2] ),
    .B1(\line_cache[138][2] ),
    .B2(_10343_),
    .X(_10908_));
 sky130_fd_sc_hd__a221o_1 _15185_ (.A1(\line_cache[137][2] ),
    .A2(_10340_),
    .B1(\line_cache[136][2] ),
    .B2(_10341_),
    .C1(_10908_),
    .X(_10909_));
 sky130_fd_sc_hd__or4_1 _15186_ (.A(_10902_),
    .B(_10905_),
    .C(_10907_),
    .D(_10909_),
    .X(_10910_));
 sky130_fd_sc_hd__nor2_1 _15187_ (.A(_10899_),
    .B(_10910_),
    .Y(_10911_));
 sky130_fd_sc_hd__and3_2 _15188_ (.A(_10860_),
    .B(_10890_),
    .C(_10911_),
    .X(_10912_));
 sky130_fd_sc_hd__and3_1 _15189_ (.A(_10772_),
    .B(_10836_),
    .C(_10912_),
    .X(_10913_));
 sky130_fd_sc_hd__nand2_1 _15190_ (.A(_09912_),
    .B(\line_cache[0][2] ),
    .Y(_10914_));
 sky130_fd_sc_hd__a21oi_4 _15191_ (.A1(_10913_),
    .A2(_10914_),
    .B1(_08979_),
    .Y(net128));
 sky130_fd_sc_hd__and2_1 _15192_ (.A(_09912_),
    .B(\line_cache[0][3] ),
    .X(_10915_));
 sky130_fd_sc_hd__and3_1 _15193_ (.A(_10102_),
    .B(\line_cache[70][3] ),
    .C(_10161_),
    .X(_10916_));
 sky130_fd_sc_hd__a22o_1 _15194_ (.A1(_10163_),
    .A2(\line_cache[68][3] ),
    .B1(_10164_),
    .B2(\line_cache[69][3] ),
    .X(_10917_));
 sky130_fd_sc_hd__a211o_1 _15195_ (.A1(\line_cache[71][3] ),
    .A2(_10159_),
    .B1(_10916_),
    .C1(_10917_),
    .X(_10918_));
 sky130_fd_sc_hd__and3_1 _15196_ (.A(_10031_),
    .B(\line_cache[77][3] ),
    .C(_10167_),
    .X(_10919_));
 sky130_fd_sc_hd__and3_1 _15197_ (.A(_10038_),
    .B(\line_cache[78][3] ),
    .C(_10167_),
    .X(_10920_));
 sky130_fd_sc_hd__and3_1 _15198_ (.A(_10041_),
    .B(\line_cache[76][3] ),
    .C(_10161_),
    .X(_10921_));
 sky130_fd_sc_hd__a2111o_1 _15199_ (.A1(_10168_),
    .A2(\line_cache[79][3] ),
    .B1(_10919_),
    .C1(_10920_),
    .D1(_10921_),
    .X(_10922_));
 sky130_fd_sc_hd__and3_1 _15200_ (.A(_10176_),
    .B(\line_cache[73][3] ),
    .C(_10167_),
    .X(_10923_));
 sky130_fd_sc_hd__a21o_1 _15201_ (.A1(\line_cache[72][3] ),
    .A2(_10175_),
    .B1(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__a221o_1 _15202_ (.A1(\line_cache[75][3] ),
    .A2(_10173_),
    .B1(\line_cache[74][3] ),
    .B2(_10174_),
    .C1(_10924_),
    .X(_10925_));
 sky130_fd_sc_hd__a22o_1 _15203_ (.A1(_10182_),
    .A2(\line_cache[64][3] ),
    .B1(_10183_),
    .B2(\line_cache[65][3] ),
    .X(_10926_));
 sky130_fd_sc_hd__a221o_1 _15204_ (.A1(\line_cache[67][3] ),
    .A2(_10180_),
    .B1(\line_cache[66][3] ),
    .B2(_10181_),
    .C1(_10926_),
    .X(_10927_));
 sky130_fd_sc_hd__or4_2 _15205_ (.A(_10918_),
    .B(_10922_),
    .C(_10925_),
    .D(_10927_),
    .X(_10928_));
 sky130_fd_sc_hd__a22o_1 _15206_ (.A1(_10189_),
    .A2(\line_cache[252][3] ),
    .B1(_10190_),
    .B2(\line_cache[251][3] ),
    .X(_10929_));
 sky130_fd_sc_hd__a221o_1 _15207_ (.A1(\line_cache[254][3] ),
    .A2(_10187_),
    .B1(\line_cache[253][3] ),
    .B2(_10188_),
    .C1(_10929_),
    .X(_10930_));
 sky130_fd_sc_hd__a22o_1 _15208_ (.A1(_10195_),
    .A2(\line_cache[248][3] ),
    .B1(_10196_),
    .B2(\line_cache[247][3] ),
    .X(_10931_));
 sky130_fd_sc_hd__a221o_1 _15209_ (.A1(\line_cache[250][3] ),
    .A2(_10193_),
    .B1(\line_cache[249][3] ),
    .B2(_10194_),
    .C1(_10931_),
    .X(_10932_));
 sky130_fd_sc_hd__and2b_1 _15210_ (.A_N(_10200_),
    .B(\line_cache[240][3] ),
    .X(_10933_));
 sky130_fd_sc_hd__and2b_1 _15211_ (.A_N(_09570_),
    .B(\line_cache[241][3] ),
    .X(_10934_));
 sky130_fd_sc_hd__and2b_1 _15212_ (.A_N(_10203_),
    .B(\line_cache[242][3] ),
    .X(_10935_));
 sky130_fd_sc_hd__a2111o_1 _15213_ (.A1(\line_cache[239][3] ),
    .A2(_10199_),
    .B1(_10933_),
    .C1(_10934_),
    .D1(_10935_),
    .X(_10936_));
 sky130_fd_sc_hd__and2b_1 _15214_ (.A_N(_10206_),
    .B(\line_cache[243][3] ),
    .X(_10937_));
 sky130_fd_sc_hd__and2b_1 _15215_ (.A_N(_10208_),
    .B(\line_cache[244][3] ),
    .X(_10938_));
 sky130_fd_sc_hd__and2b_1 _15216_ (.A_N(_09597_),
    .B(\line_cache[245][3] ),
    .X(_10939_));
 sky130_fd_sc_hd__and2b_1 _15217_ (.A_N(_10211_),
    .B(\line_cache[246][3] ),
    .X(_10940_));
 sky130_fd_sc_hd__or4_1 _15218_ (.A(_10937_),
    .B(_10938_),
    .C(_10939_),
    .D(_10940_),
    .X(_10941_));
 sky130_fd_sc_hd__or4_1 _15219_ (.A(_10930_),
    .B(_10932_),
    .C(_10936_),
    .D(_10941_),
    .X(_10942_));
 sky130_fd_sc_hd__and3_1 _15220_ (.A(_09595_),
    .B(\line_cache[229][3] ),
    .C(_10099_),
    .X(_10943_));
 sky130_fd_sc_hd__and3_1 _15221_ (.A(_10102_),
    .B(\line_cache[230][3] ),
    .C(_10434_),
    .X(_10944_));
 sky130_fd_sc_hd__and3_1 _15222_ (.A(_10104_),
    .B(\line_cache[227][3] ),
    .C(_10434_),
    .X(_10945_));
 sky130_fd_sc_hd__and3_1 _15223_ (.A(_10106_),
    .B(\line_cache[228][3] ),
    .C(_10437_),
    .X(_10946_));
 sky130_fd_sc_hd__or4_1 _15224_ (.A(_10943_),
    .B(_10944_),
    .C(_10945_),
    .D(_10946_),
    .X(_10947_));
 sky130_fd_sc_hd__and3_1 _15225_ (.A(_09544_),
    .B(\line_cache[223][3] ),
    .C(_10109_),
    .X(_10948_));
 sky130_fd_sc_hd__and3_1 _15226_ (.A(_10071_),
    .B(\line_cache[224][3] ),
    .C(_10434_),
    .X(_10949_));
 sky130_fd_sc_hd__and3_1 _15227_ (.A(_10067_),
    .B(\line_cache[225][3] ),
    .C(_10437_),
    .X(_10950_));
 sky130_fd_sc_hd__and3_1 _15228_ (.A(_10074_),
    .B(\line_cache[226][3] ),
    .C(_10437_),
    .X(_10951_));
 sky130_fd_sc_hd__or4_1 _15229_ (.A(_10948_),
    .B(_10949_),
    .C(_10950_),
    .D(_10951_),
    .X(_10952_));
 sky130_fd_sc_hd__a22o_1 _15230_ (.A1(_10118_),
    .A2(\line_cache[236][3] ),
    .B1(_10120_),
    .B2(\line_cache[235][3] ),
    .X(_10953_));
 sky130_fd_sc_hd__a221o_1 _15231_ (.A1(\line_cache[238][3] ),
    .A2(_10116_),
    .B1(\line_cache[237][3] ),
    .B2(_10117_),
    .C1(_10953_),
    .X(_10954_));
 sky130_fd_sc_hd__a22o_1 _15232_ (.A1(_10125_),
    .A2(\line_cache[232][3] ),
    .B1(_10126_),
    .B2(\line_cache[231][3] ),
    .X(_10955_));
 sky130_fd_sc_hd__a221o_1 _15233_ (.A1(\line_cache[234][3] ),
    .A2(_10123_),
    .B1(\line_cache[233][3] ),
    .B2(_10124_),
    .C1(_10955_),
    .X(_10956_));
 sky130_fd_sc_hd__or4_1 _15234_ (.A(_10947_),
    .B(_10952_),
    .C(_10954_),
    .D(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__a22o_1 _15235_ (.A1(_10132_),
    .A2(\line_cache[220][3] ),
    .B1(_10133_),
    .B2(\line_cache[219][3] ),
    .X(_10958_));
 sky130_fd_sc_hd__a221o_1 _15236_ (.A1(\line_cache[222][3] ),
    .A2(_10130_),
    .B1(\line_cache[221][3] ),
    .B2(_10131_),
    .C1(_10958_),
    .X(_10959_));
 sky130_fd_sc_hd__a22o_1 _15237_ (.A1(_10138_),
    .A2(\line_cache[208][3] ),
    .B1(_10139_),
    .B2(\line_cache[207][3] ),
    .X(_10960_));
 sky130_fd_sc_hd__a221o_1 _15238_ (.A1(\line_cache[210][3] ),
    .A2(_10136_),
    .B1(\line_cache[209][3] ),
    .B2(_10137_),
    .C1(_10960_),
    .X(_10961_));
 sky130_fd_sc_hd__a22o_1 _15239_ (.A1(_10144_),
    .A2(\line_cache[216][3] ),
    .B1(_10145_),
    .B2(\line_cache[215][3] ),
    .X(_10962_));
 sky130_fd_sc_hd__a221o_1 _15240_ (.A1(\line_cache[218][3] ),
    .A2(_10142_),
    .B1(\line_cache[217][3] ),
    .B2(_10143_),
    .C1(_10962_),
    .X(_10963_));
 sky130_fd_sc_hd__and2b_1 _15241_ (.A_N(_10148_),
    .B(\line_cache[211][3] ),
    .X(_10964_));
 sky130_fd_sc_hd__nor2b_1 _15242_ (.A(_10150_),
    .B_N(\line_cache[212][3] ),
    .Y(_10965_));
 sky130_fd_sc_hd__and2b_1 _15243_ (.A_N(_10152_),
    .B(\line_cache[213][3] ),
    .X(_10966_));
 sky130_fd_sc_hd__and2b_1 _15244_ (.A_N(_10154_),
    .B(\line_cache[214][3] ),
    .X(_10967_));
 sky130_fd_sc_hd__or4_1 _15245_ (.A(_10964_),
    .B(_10965_),
    .C(_10966_),
    .D(_10967_),
    .X(_10968_));
 sky130_fd_sc_hd__or4_1 _15246_ (.A(_10959_),
    .B(_10961_),
    .C(_10963_),
    .D(_10968_),
    .X(_10969_));
 sky130_fd_sc_hd__or2_1 _15247_ (.A(_10957_),
    .B(_10969_),
    .X(_10970_));
 sky130_fd_sc_hd__or3_2 _15248_ (.A(_10928_),
    .B(_10942_),
    .C(_10970_),
    .X(_10971_));
 sky130_fd_sc_hd__and3_1 _15249_ (.A(_10035_),
    .B(\line_cache[203][3] ),
    .C(_09539_),
    .X(_10972_));
 sky130_fd_sc_hd__and3_1 _15250_ (.A(_10038_),
    .B(\line_cache[206][3] ),
    .C(_10075_),
    .X(_10973_));
 sky130_fd_sc_hd__and3_1 _15251_ (.A(_10041_),
    .B(\line_cache[204][3] ),
    .C(_10075_),
    .X(_10974_));
 sky130_fd_sc_hd__a2111o_1 _15252_ (.A1(\line_cache[205][3] ),
    .A2(_10033_),
    .B1(_10972_),
    .C1(_10973_),
    .D1(_10974_),
    .X(_10975_));
 sky130_fd_sc_hd__a22o_1 _15253_ (.A1(_10049_),
    .A2(\line_cache[195][3] ),
    .B1(\line_cache[196][3] ),
    .B2(_10051_),
    .X(_10976_));
 sky130_fd_sc_hd__a221o_1 _15254_ (.A1(\line_cache[198][3] ),
    .A2(_10046_),
    .B1(\line_cache[197][3] ),
    .B2(_10047_),
    .C1(_10976_),
    .X(_10977_));
 sky130_fd_sc_hd__a22o_1 _15255_ (.A1(_10060_),
    .A2(\line_cache[200][3] ),
    .B1(_10063_),
    .B2(\line_cache[199][3] ),
    .X(_10978_));
 sky130_fd_sc_hd__a221o_1 _15256_ (.A1(\line_cache[202][3] ),
    .A2(_10056_),
    .B1(\line_cache[201][3] ),
    .B2(_10059_),
    .C1(_10978_),
    .X(_10979_));
 sky130_fd_sc_hd__and3_1 _15257_ (.A(_10067_),
    .B(\line_cache[193][3] ),
    .C(_09540_),
    .X(_10980_));
 sky130_fd_sc_hd__and3_1 _15258_ (.A(_10071_),
    .B(\line_cache[192][3] ),
    .C(_09540_),
    .X(_10981_));
 sky130_fd_sc_hd__and3_1 _15259_ (.A(_10074_),
    .B(\line_cache[194][3] ),
    .C(_09540_),
    .X(_10982_));
 sky130_fd_sc_hd__a2111o_1 _15260_ (.A1(_10066_),
    .A2(\line_cache[286][3] ),
    .B1(_10980_),
    .C1(_10981_),
    .D1(_10982_),
    .X(_10983_));
 sky130_fd_sc_hd__or4_1 _15261_ (.A(_10975_),
    .B(_10977_),
    .C(_10979_),
    .D(_10983_),
    .X(_10984_));
 sky130_fd_sc_hd__a22o_1 _15262_ (.A1(_09623_),
    .A2(\line_cache[275][3] ),
    .B1(_09620_),
    .B2(\line_cache[274][3] ),
    .X(_10985_));
 sky130_fd_sc_hd__a22o_1 _15263_ (.A1(_10080_),
    .A2(\line_cache[276][3] ),
    .B1(\line_cache[277][3] ),
    .B2(_10081_),
    .X(_10986_));
 sky130_fd_sc_hd__a22o_1 _15264_ (.A1(_10086_),
    .A2(\line_cache[270][3] ),
    .B1(\line_cache[269][3] ),
    .B2(_10088_),
    .X(_10987_));
 sky130_fd_sc_hd__a221o_1 _15265_ (.A1(\line_cache[273][3] ),
    .A2(_10083_),
    .B1(\line_cache[272][3] ),
    .B2(_10084_),
    .C1(_10987_),
    .X(_10988_));
 sky130_fd_sc_hd__a22o_1 _15266_ (.A1(_09658_),
    .A2(\line_cache[283][3] ),
    .B1(\line_cache[282][3] ),
    .B2(_09661_),
    .X(_10989_));
 sky130_fd_sc_hd__a22o_1 _15267_ (.A1(_09645_),
    .A2(\line_cache[285][3] ),
    .B1(\line_cache[284][3] ),
    .B2(_09648_),
    .X(_10990_));
 sky130_fd_sc_hd__a22o_1 _15268_ (.A1(_09639_),
    .A2(\line_cache[279][3] ),
    .B1(\line_cache[278][3] ),
    .B2(_09636_),
    .X(_10991_));
 sky130_fd_sc_hd__a221o_1 _15269_ (.A1(\line_cache[281][3] ),
    .A2(_09663_),
    .B1(\line_cache[280][3] ),
    .B2(_09655_),
    .C1(_10991_),
    .X(_10992_));
 sky130_fd_sc_hd__or3_1 _15270_ (.A(_10989_),
    .B(_10990_),
    .C(_10992_),
    .X(_10993_));
 sky130_fd_sc_hd__or4_1 _15271_ (.A(_10985_),
    .B(_10986_),
    .C(_10988_),
    .D(_10993_),
    .X(_10994_));
 sky130_fd_sc_hd__nor2_1 _15272_ (.A(_10984_),
    .B(_10994_),
    .Y(_10995_));
 sky130_fd_sc_hd__and2b_1 _15273_ (.A_N(_09987_),
    .B(\line_cache[256][3] ),
    .X(_10996_));
 sky130_fd_sc_hd__and2b_1 _15274_ (.A_N(_09747_),
    .B(\line_cache[302][3] ),
    .X(_10997_));
 sky130_fd_sc_hd__a22o_1 _15275_ (.A1(_09743_),
    .A2(\line_cache[301][3] ),
    .B1(\line_cache[300][3] ),
    .B2(_09742_),
    .X(_10998_));
 sky130_fd_sc_hd__or3_1 _15276_ (.A(_10996_),
    .B(_10997_),
    .C(_10998_),
    .X(_10999_));
 sky130_fd_sc_hd__and3_1 _15277_ (.A(_09917_),
    .B(_09691_),
    .C(\line_cache[258][3] ),
    .X(_11000_));
 sky130_fd_sc_hd__and3_1 _15278_ (.A(_09848_),
    .B(_09691_),
    .C(\line_cache[260][3] ),
    .X(_11001_));
 sky130_fd_sc_hd__and3_1 _15279_ (.A(_09919_),
    .B(_09611_),
    .C(\line_cache[257][3] ),
    .X(_11002_));
 sky130_fd_sc_hd__and3_1 _15280_ (.A(_09840_),
    .B(_09611_),
    .C(\line_cache[259][3] ),
    .X(_11003_));
 sky130_fd_sc_hd__or4_1 _15281_ (.A(_11000_),
    .B(_11001_),
    .C(_11002_),
    .D(_11003_),
    .X(_11004_));
 sky130_fd_sc_hd__and3_1 _15282_ (.A(_09858_),
    .B(_09547_),
    .C(\line_cache[267][3] ),
    .X(_11005_));
 sky130_fd_sc_hd__a22o_1 _15283_ (.A1(_09998_),
    .A2(\line_cache[265][3] ),
    .B1(\line_cache[266][3] ),
    .B2(_09999_),
    .X(_11006_));
 sky130_fd_sc_hd__a311o_1 _15284_ (.A1(_09548_),
    .A2(\line_cache[268][3] ),
    .A3(_09862_),
    .B1(_11005_),
    .C1(_11006_),
    .X(_11007_));
 sky130_fd_sc_hd__nand2_1 _15285_ (.A(_10007_),
    .B(\line_cache[262][3] ),
    .Y(_11008_));
 sky130_fd_sc_hd__nand2_1 _15286_ (.A(_10010_),
    .B(\line_cache[261][3] ),
    .Y(_11009_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(_11008_),
    .B(_11009_),
    .Y(_11010_));
 sky130_fd_sc_hd__a221oi_1 _15288_ (.A1(_10003_),
    .A2(\line_cache[264][3] ),
    .B1(_10005_),
    .B2(\line_cache[263][3] ),
    .C1(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__or4b_1 _15289_ (.A(_10999_),
    .B(_11004_),
    .C(_11007_),
    .D_N(_11011_),
    .X(_11012_));
 sky130_fd_sc_hd__a22o_1 _15290_ (.A1(_09682_),
    .A2(\line_cache[308][3] ),
    .B1(\line_cache[309][3] ),
    .B2(_09685_),
    .X(_11013_));
 sky130_fd_sc_hd__a221o_1 _15291_ (.A1(\line_cache[311][3] ),
    .A2(_09689_),
    .B1(\line_cache[310][3] ),
    .B2(_09693_),
    .C1(_11013_),
    .X(_11014_));
 sky130_fd_sc_hd__a22o_1 _15292_ (.A1(_09728_),
    .A2(\line_cache[295][3] ),
    .B1(\line_cache[294][3] ),
    .B2(_09726_),
    .X(_11015_));
 sky130_fd_sc_hd__a221o_1 _15293_ (.A1(\line_cache[293][3] ),
    .A2(_09730_),
    .B1(\line_cache[292][3] ),
    .B2(_10018_),
    .C1(_11015_),
    .X(_11016_));
 sky130_fd_sc_hd__a22o_1 _15294_ (.A1(_09716_),
    .A2(\line_cache[296][3] ),
    .B1(\line_cache[297][3] ),
    .B2(_09721_),
    .X(_11017_));
 sky130_fd_sc_hd__a221o_1 _15295_ (.A1(\line_cache[299][3] ),
    .A2(_09718_),
    .B1(\line_cache[298][3] ),
    .B2(_09720_),
    .C1(_11017_),
    .X(_11018_));
 sky130_fd_sc_hd__a22o_1 _15296_ (.A1(_10025_),
    .A2(\line_cache[288][3] ),
    .B1(\line_cache[289][3] ),
    .B2(_10026_),
    .X(_11019_));
 sky130_fd_sc_hd__a221o_1 _15297_ (.A1(\line_cache[291][3] ),
    .A2(_10023_),
    .B1(\line_cache[290][3] ),
    .B2(_10024_),
    .C1(_11019_),
    .X(_11020_));
 sky130_fd_sc_hd__or4_4 _15298_ (.A(_11014_),
    .B(_11016_),
    .C(_11018_),
    .D(_11020_),
    .X(_11021_));
 sky130_fd_sc_hd__nor2_1 _15299_ (.A(_11012_),
    .B(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__nand2_1 _15300_ (.A(_10995_),
    .B(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__nor2_1 _15301_ (.A(_10971_),
    .B(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__a22o_1 _15302_ (.A1(_09842_),
    .A2(\line_cache[6][3] ),
    .B1(\line_cache[5][3] ),
    .B2(_09844_),
    .X(_11025_));
 sky130_fd_sc_hd__a221o_1 _15303_ (.A1(\line_cache[4][3] ),
    .A2(_09850_),
    .B1(\line_cache[3][3] ),
    .B2(_09914_),
    .C1(_11025_),
    .X(_11026_));
 sky130_fd_sc_hd__and3_1 _15304_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][3] ),
    .X(_11027_));
 sky130_fd_sc_hd__and3_1 _15305_ (.A(_09919_),
    .B(_09533_),
    .C(\line_cache[1][3] ),
    .X(_11028_));
 sky130_fd_sc_hd__a211o_1 _15306_ (.A1(\line_cache[15][3] ),
    .A2(_09867_),
    .B1(_11027_),
    .C1(_11028_),
    .X(_11029_));
 sky130_fd_sc_hd__and3_1 _15307_ (.A(_09922_),
    .B(_09532_),
    .C(\line_cache[63][3] ),
    .X(_11030_));
 sky130_fd_sc_hd__a31o_1 _15308_ (.A1(_09548_),
    .A2(\line_cache[319][3] ),
    .A3(_09922_),
    .B1(_11030_),
    .X(_11031_));
 sky130_fd_sc_hd__a221o_1 _15309_ (.A1(\line_cache[47][3] ),
    .A2(_09806_),
    .B1(\line_cache[31][3] ),
    .B2(_09907_),
    .C1(_11031_),
    .X(_11032_));
 sky130_fd_sc_hd__nand2_1 _15310_ (.A(_09746_),
    .B(\line_cache[303][3] ),
    .Y(_11033_));
 sky130_fd_sc_hd__nand2_1 _15311_ (.A(_09930_),
    .B(\line_cache[271][3] ),
    .Y(_11034_));
 sky130_fd_sc_hd__nand2_1 _15312_ (.A(_11033_),
    .B(_11034_),
    .Y(_11035_));
 sky130_fd_sc_hd__a221oi_2 _15313_ (.A1(\line_cache[255][3] ),
    .A2(_09926_),
    .B1(\line_cache[287][3] ),
    .B2(_09927_),
    .C1(_11035_),
    .Y(_11036_));
 sky130_fd_sc_hd__or4b_1 _15314_ (.A(_11026_),
    .B(_11029_),
    .C(_11032_),
    .D_N(_11036_),
    .X(_11037_));
 sky130_fd_sc_hd__a22o_1 _15315_ (.A1(_09803_),
    .A2(\line_cache[45][3] ),
    .B1(\line_cache[46][3] ),
    .B2(_09804_),
    .X(_11038_));
 sky130_fd_sc_hd__a22o_1 _15316_ (.A1(_09824_),
    .A2(\line_cache[48][3] ),
    .B1(\line_cache[49][3] ),
    .B2(_09826_),
    .X(_11039_));
 sky130_fd_sc_hd__nand2_1 _15317_ (.A(_09787_),
    .B(\line_cache[41][3] ),
    .Y(_11040_));
 sky130_fd_sc_hd__nand2_1 _15318_ (.A(_09789_),
    .B(\line_cache[42][3] ),
    .Y(_11041_));
 sky130_fd_sc_hd__nand2_1 _15319_ (.A(_11040_),
    .B(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__a221oi_2 _15320_ (.A1(_09785_),
    .A2(\line_cache[43][3] ),
    .B1(\line_cache[44][3] ),
    .B2(_09801_),
    .C1(_11042_),
    .Y(_11043_));
 sky130_fd_sc_hd__or3b_1 _15321_ (.A(_11038_),
    .B(_11039_),
    .C_N(_11043_),
    .X(_11044_));
 sky130_fd_sc_hd__a22o_1 _15322_ (.A1(_09699_),
    .A2(\line_cache[317][3] ),
    .B1(\line_cache[316][3] ),
    .B2(_09697_),
    .X(_11045_));
 sky130_fd_sc_hd__a22o_1 _15323_ (.A1(_09832_),
    .A2(\line_cache[58][3] ),
    .B1(\line_cache[59][3] ),
    .B2(_09833_),
    .X(_11046_));
 sky130_fd_sc_hd__a22o_1 _15324_ (.A1(_09819_),
    .A2(\line_cache[61][3] ),
    .B1(\line_cache[60][3] ),
    .B2(_09817_),
    .X(_11047_));
 sky130_fd_sc_hd__a22o_1 _15325_ (.A1(_09822_),
    .A2(\line_cache[62][3] ),
    .B1(\line_cache[318][3] ),
    .B2(_09702_),
    .X(_11048_));
 sky130_fd_sc_hd__or4_2 _15326_ (.A(_11045_),
    .B(_11046_),
    .C(_11047_),
    .D(_11048_),
    .X(_11049_));
 sky130_fd_sc_hd__a22o_1 _15327_ (.A1(_09675_),
    .A2(\line_cache[304][3] ),
    .B1(\line_cache[305][3] ),
    .B2(_09676_),
    .X(_11050_));
 sky130_fd_sc_hd__a22o_1 _15328_ (.A1(_09705_),
    .A2(\line_cache[312][3] ),
    .B1(\line_cache[313][3] ),
    .B2(_09707_),
    .X(_11051_));
 sky130_fd_sc_hd__a22o_1 _15329_ (.A1(_09708_),
    .A2(\line_cache[314][3] ),
    .B1(\line_cache[315][3] ),
    .B2(_09709_),
    .X(_11052_));
 sky130_fd_sc_hd__a22o_1 _15330_ (.A1(_09677_),
    .A2(\line_cache[306][3] ),
    .B1(\line_cache[307][3] ),
    .B2(_09678_),
    .X(_11053_));
 sky130_fd_sc_hd__or4_1 _15331_ (.A(_11050_),
    .B(_11051_),
    .C(_11052_),
    .D(_11053_),
    .X(_11054_));
 sky130_fd_sc_hd__a22o_1 _15332_ (.A1(_09830_),
    .A2(\line_cache[56][3] ),
    .B1(\line_cache[57][3] ),
    .B2(_09834_),
    .X(_11055_));
 sky130_fd_sc_hd__a22o_1 _15333_ (.A1(_09809_),
    .A2(\line_cache[52][3] ),
    .B1(\line_cache[53][3] ),
    .B2(_09811_),
    .X(_11056_));
 sky130_fd_sc_hd__a22o_1 _15334_ (.A1(_09827_),
    .A2(\line_cache[50][3] ),
    .B1(\line_cache[51][3] ),
    .B2(_09828_),
    .X(_11057_));
 sky130_fd_sc_hd__a22o_1 _15335_ (.A1(_09813_),
    .A2(\line_cache[54][3] ),
    .B1(\line_cache[55][3] ),
    .B2(_09815_),
    .X(_11058_));
 sky130_fd_sc_hd__or4_1 _15336_ (.A(_11055_),
    .B(_11056_),
    .C(_11057_),
    .D(_11058_),
    .X(_11059_));
 sky130_fd_sc_hd__or4_2 _15337_ (.A(_11044_),
    .B(_11049_),
    .C(_11054_),
    .D(_11059_),
    .X(_11060_));
 sky130_fd_sc_hd__nand2_1 _15338_ (.A(_09864_),
    .B(\line_cache[12][3] ),
    .Y(_11061_));
 sky130_fd_sc_hd__nand2_1 _15339_ (.A(_09860_),
    .B(\line_cache[11][3] ),
    .Y(_11062_));
 sky130_fd_sc_hd__nand2_1 _15340_ (.A(_11061_),
    .B(_11062_),
    .Y(_11063_));
 sky130_fd_sc_hd__a221oi_1 _15341_ (.A1(_09870_),
    .A2(\line_cache[14][3] ),
    .B1(\line_cache[13][3] ),
    .B2(_09873_),
    .C1(_11063_),
    .Y(_11064_));
 sky130_fd_sc_hd__nand2_1 _15342_ (.A(_09853_),
    .B(\line_cache[10][3] ),
    .Y(_11065_));
 sky130_fd_sc_hd__nand2_1 _15343_ (.A(_09857_),
    .B(\line_cache[9][3] ),
    .Y(_11066_));
 sky130_fd_sc_hd__nand2_1 _15344_ (.A(_11065_),
    .B(_11066_),
    .Y(_11067_));
 sky130_fd_sc_hd__a221oi_1 _15345_ (.A1(_09855_),
    .A2(\line_cache[8][3] ),
    .B1(_09847_),
    .B2(\line_cache[7][3] ),
    .C1(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__nand2_1 _15346_ (.A(_11064_),
    .B(_11068_),
    .Y(_11069_));
 sky130_fd_sc_hd__and3_1 _15347_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][3] ),
    .X(_11070_));
 sky130_fd_sc_hd__a22o_1 _15348_ (.A1(_09884_),
    .A2(\line_cache[23][3] ),
    .B1(\line_cache[22][3] ),
    .B2(_09886_),
    .X(_11071_));
 sky130_fd_sc_hd__a22o_1 _15349_ (.A1(_09877_),
    .A2(\line_cache[19][3] ),
    .B1(\line_cache[18][3] ),
    .B2(_09878_),
    .X(_11072_));
 sky130_fd_sc_hd__a221o_1 _15350_ (.A1(\line_cache[17][3] ),
    .A2(_09969_),
    .B1(\line_cache[16][3] ),
    .B2(_09970_),
    .C1(_11072_),
    .X(_11073_));
 sky130_fd_sc_hd__a2111o_1 _15351_ (.A1(\line_cache[20][3] ),
    .A2(_09888_),
    .B1(_11070_),
    .C1(_11071_),
    .D1(_11073_),
    .X(_11074_));
 sky130_fd_sc_hd__a22o_1 _15352_ (.A1(_09796_),
    .A2(\line_cache[33][3] ),
    .B1(\line_cache[34][3] ),
    .B2(_09798_),
    .X(_11075_));
 sky130_fd_sc_hd__a221o_1 _15353_ (.A1(\line_cache[36][3] ),
    .A2(_09777_),
    .B1(\line_cache[35][3] ),
    .B2(_09794_),
    .C1(_11075_),
    .X(_11076_));
 sky130_fd_sc_hd__a22o_1 _15354_ (.A1(_09890_),
    .A2(\line_cache[27][3] ),
    .B1(\line_cache[26][3] ),
    .B2(_09896_),
    .X(_11077_));
 sky130_fd_sc_hd__a221oi_2 _15355_ (.A1(\line_cache[25][3] ),
    .A2(_09892_),
    .B1(\line_cache[24][3] ),
    .B2(_09895_),
    .C1(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__a22o_1 _15356_ (.A1(_09903_),
    .A2(\line_cache[29][3] ),
    .B1(\line_cache[28][3] ),
    .B2(_09900_),
    .X(_11079_));
 sky130_fd_sc_hd__a221oi_1 _15357_ (.A1(\line_cache[32][3] ),
    .A2(_09792_),
    .B1(\line_cache[30][3] ),
    .B2(_09905_),
    .C1(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__nand2_1 _15358_ (.A(_09773_),
    .B(\line_cache[38][3] ),
    .Y(_11081_));
 sky130_fd_sc_hd__nand2_1 _15359_ (.A(_09775_),
    .B(\line_cache[37][3] ),
    .Y(_11082_));
 sky130_fd_sc_hd__nand2_1 _15360_ (.A(_11081_),
    .B(_11082_),
    .Y(_11083_));
 sky130_fd_sc_hd__a221oi_2 _15361_ (.A1(_09783_),
    .A2(\line_cache[40][3] ),
    .B1(\line_cache[39][3] ),
    .B2(_09780_),
    .C1(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__and4b_1 _15362_ (.A_N(_11076_),
    .B(_11078_),
    .C(_11080_),
    .D(_11084_),
    .X(_11085_));
 sky130_fd_sc_hd__or3b_1 _15363_ (.A(_11069_),
    .B(_11074_),
    .C_N(_11085_),
    .X(_11086_));
 sky130_fd_sc_hd__nor3_1 _15364_ (.A(_11037_),
    .B(_11060_),
    .C(_11086_),
    .Y(_11087_));
 sky130_fd_sc_hd__a22o_1 _15365_ (.A1(_10244_),
    .A2(\line_cache[173][3] ),
    .B1(\line_cache[172][3] ),
    .B2(_10245_),
    .X(_11088_));
 sky130_fd_sc_hd__a221o_1 _15366_ (.A1(\line_cache[175][3] ),
    .A2(_10242_),
    .B1(\line_cache[174][3] ),
    .B2(_10243_),
    .C1(_11088_),
    .X(_11089_));
 sky130_fd_sc_hd__a22o_1 _15367_ (.A1(_10263_),
    .A2(\line_cache[170][3] ),
    .B1(\line_cache[171][3] ),
    .B2(_10262_),
    .X(_11090_));
 sky130_fd_sc_hd__a221o_1 _15368_ (.A1(\line_cache[169][3] ),
    .A2(_10260_),
    .B1(\line_cache[168][3] ),
    .B2(_10261_),
    .C1(_11090_),
    .X(_11091_));
 sky130_fd_sc_hd__a22o_1 _15369_ (.A1(_10256_),
    .A2(\line_cache[160][3] ),
    .B1(\line_cache[161][3] ),
    .B2(_10257_),
    .X(_11092_));
 sky130_fd_sc_hd__and3_1 _15370_ (.A(_10104_),
    .B(_09751_),
    .C(\line_cache[163][3] ),
    .X(_11093_));
 sky130_fd_sc_hd__a22o_1 _15371_ (.A1(_10249_),
    .A2(\line_cache[166][3] ),
    .B1(\line_cache[167][3] ),
    .B2(_10248_),
    .X(_11094_));
 sky130_fd_sc_hd__a221o_1 _15372_ (.A1(\line_cache[165][3] ),
    .A2(_10250_),
    .B1(\line_cache[164][3] ),
    .B2(_10251_),
    .C1(_11094_),
    .X(_11095_));
 sky130_fd_sc_hd__a2111o_1 _15373_ (.A1(\line_cache[162][3] ),
    .A2(_10255_),
    .B1(_11092_),
    .C1(_11093_),
    .D1(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__nor3_1 _15374_ (.A(_11089_),
    .B(_11091_),
    .C(_11096_),
    .Y(_11097_));
 sky130_fd_sc_hd__a22o_1 _15375_ (.A1(_10277_),
    .A2(\line_cache[184][3] ),
    .B1(\line_cache[185][3] ),
    .B2(_10278_),
    .X(_11098_));
 sky130_fd_sc_hd__a221o_1 _15376_ (.A1(\line_cache[187][3] ),
    .A2(_10275_),
    .B1(\line_cache[186][3] ),
    .B2(_10276_),
    .C1(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__a22o_1 _15377_ (.A1(_10284_),
    .A2(\line_cache[176][3] ),
    .B1(_10285_),
    .B2(\line_cache[177][3] ),
    .X(_11100_));
 sky130_fd_sc_hd__a221oi_1 _15378_ (.A1(\line_cache[179][3] ),
    .A2(_10282_),
    .B1(\line_cache[178][3] ),
    .B2(_10283_),
    .C1(_11100_),
    .Y(_11101_));
 sky130_fd_sc_hd__and3_1 _15379_ (.A(_10288_),
    .B(_10102_),
    .C(\line_cache[182][3] ),
    .X(_11102_));
 sky130_fd_sc_hd__and3_1 _15380_ (.A(_10288_),
    .B(_10098_),
    .C(\line_cache[181][3] ),
    .X(_11103_));
 sky130_fd_sc_hd__a31o_1 _15381_ (.A1(\line_cache[180][3] ),
    .A2(_10289_),
    .A3(_10106_),
    .B1(_11103_),
    .X(_11104_));
 sky130_fd_sc_hd__a311oi_2 _15382_ (.A1(\line_cache[183][3] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_11102_),
    .C1(_11104_),
    .Y(_11105_));
 sky130_fd_sc_hd__a22o_1 _15383_ (.A1(_10272_),
    .A2(\line_cache[189][3] ),
    .B1(\line_cache[188][3] ),
    .B2(_10271_),
    .X(_11106_));
 sky130_fd_sc_hd__a221oi_1 _15384_ (.A1(\line_cache[191][3] ),
    .A2(_10269_),
    .B1(\line_cache[190][3] ),
    .B2(_10270_),
    .C1(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__and4b_1 _15385_ (.A_N(_11099_),
    .B(_11101_),
    .C(_11105_),
    .D(_11107_),
    .X(_11108_));
 sky130_fd_sc_hd__a22o_1 _15386_ (.A1(_10219_),
    .A2(\line_cache[157][3] ),
    .B1(\line_cache[156][3] ),
    .B2(_10220_),
    .X(_11109_));
 sky130_fd_sc_hd__a221o_1 _15387_ (.A1(\line_cache[159][3] ),
    .A2(_10217_),
    .B1(\line_cache[158][3] ),
    .B2(_10218_),
    .C1(_11109_),
    .X(_11110_));
 sky130_fd_sc_hd__a22o_1 _15388_ (.A1(_10238_),
    .A2(\line_cache[154][3] ),
    .B1(\line_cache[155][3] ),
    .B2(_10237_),
    .X(_11111_));
 sky130_fd_sc_hd__a221o_1 _15389_ (.A1(\line_cache[153][3] ),
    .A2(_10235_),
    .B1(\line_cache[152][3] ),
    .B2(_10236_),
    .C1(_11111_),
    .X(_11112_));
 sky130_fd_sc_hd__a22o_1 _15390_ (.A1(_10224_),
    .A2(\line_cache[148][3] ),
    .B1(\line_cache[149][3] ),
    .B2(_10223_),
    .X(_11113_));
 sky130_fd_sc_hd__a22o_1 _15391_ (.A1(_10225_),
    .A2(\line_cache[151][3] ),
    .B1(\line_cache[150][3] ),
    .B2(_10226_),
    .X(_11114_));
 sky130_fd_sc_hd__a22o_1 _15392_ (.A1(_10230_),
    .A2(\line_cache[144][3] ),
    .B1(\line_cache[145][3] ),
    .B2(_10229_),
    .X(_11115_));
 sky130_fd_sc_hd__a22o_1 _15393_ (.A1(_10231_),
    .A2(\line_cache[147][3] ),
    .B1(\line_cache[146][3] ),
    .B2(_10232_),
    .X(_11116_));
 sky130_fd_sc_hd__or4_1 _15394_ (.A(_11113_),
    .B(_11114_),
    .C(_11115_),
    .D(_11116_),
    .X(_11117_));
 sky130_fd_sc_hd__nor3_1 _15395_ (.A(_11110_),
    .B(_11112_),
    .C(_11117_),
    .Y(_11118_));
 sky130_fd_sc_hd__and3_2 _15396_ (.A(_11097_),
    .B(_11108_),
    .C(_11118_),
    .X(_11119_));
 sky130_fd_sc_hd__a22o_1 _15397_ (.A1(_10378_),
    .A2(\line_cache[80][3] ),
    .B1(_10379_),
    .B2(\line_cache[81][3] ),
    .X(_11120_));
 sky130_fd_sc_hd__a221o_1 _15398_ (.A1(\line_cache[83][3] ),
    .A2(_10376_),
    .B1(\line_cache[82][3] ),
    .B2(_10377_),
    .C1(_11120_),
    .X(_11121_));
 sky130_fd_sc_hd__a22o_1 _15399_ (.A1(_10384_),
    .A2(\line_cache[92][3] ),
    .B1(_10385_),
    .B2(\line_cache[93][3] ),
    .X(_11122_));
 sky130_fd_sc_hd__a221o_1 _15400_ (.A1(\line_cache[95][3] ),
    .A2(net136),
    .B1(\line_cache[94][3] ),
    .B2(_10383_),
    .C1(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__a22o_1 _15401_ (.A1(_10390_),
    .A2(\line_cache[84][3] ),
    .B1(_10391_),
    .B2(\line_cache[85][3] ),
    .X(_11124_));
 sky130_fd_sc_hd__a221o_1 _15402_ (.A1(\line_cache[87][3] ),
    .A2(_10388_),
    .B1(\line_cache[86][3] ),
    .B2(_10389_),
    .C1(_11124_),
    .X(_11125_));
 sky130_fd_sc_hd__a22o_1 _15403_ (.A1(_10396_),
    .A2(\line_cache[88][3] ),
    .B1(_10397_),
    .B2(\line_cache[89][3] ),
    .X(_11126_));
 sky130_fd_sc_hd__a221o_1 _15404_ (.A1(\line_cache[91][3] ),
    .A2(_10394_),
    .B1(\line_cache[90][3] ),
    .B2(_10395_),
    .C1(_11126_),
    .X(_11127_));
 sky130_fd_sc_hd__or4_1 _15405_ (.A(_11121_),
    .B(_11123_),
    .C(_11125_),
    .D(_11127_),
    .X(_11128_));
 sky130_fd_sc_hd__a22o_1 _15406_ (.A1(_10371_),
    .A2(\line_cache[100][3] ),
    .B1(_10372_),
    .B2(\line_cache[101][3] ),
    .X(_11129_));
 sky130_fd_sc_hd__a22o_1 _15407_ (.A1(_10369_),
    .A2(\line_cache[103][3] ),
    .B1(_10370_),
    .B2(\line_cache[102][3] ),
    .X(_11130_));
 sky130_fd_sc_hd__a22o_1 _15408_ (.A1(_10351_),
    .A2(\line_cache[96][3] ),
    .B1(_10352_),
    .B2(\line_cache[97][3] ),
    .X(_11131_));
 sky130_fd_sc_hd__a221o_2 _15409_ (.A1(\line_cache[99][3] ),
    .A2(_10349_),
    .B1(\line_cache[98][3] ),
    .B2(_10348_),
    .C1(_11131_),
    .X(_11132_));
 sky130_fd_sc_hd__and3_1 _15410_ (.A(_10035_),
    .B(\line_cache[107][3] ),
    .C(_10651_),
    .X(_11133_));
 sky130_fd_sc_hd__and3_1 _15411_ (.A(_10176_),
    .B(\line_cache[105][3] ),
    .C(_10651_),
    .X(_11134_));
 sky130_fd_sc_hd__and3_1 _15412_ (.A(_10054_),
    .B(\line_cache[106][3] ),
    .C(_10356_),
    .X(_11135_));
 sky130_fd_sc_hd__and3_1 _15413_ (.A(_10360_),
    .B(\line_cache[104][3] ),
    .C(_10356_),
    .X(_11136_));
 sky130_fd_sc_hd__or4_1 _15414_ (.A(_11133_),
    .B(_11134_),
    .C(_11135_),
    .D(_11136_),
    .X(_11137_));
 sky130_fd_sc_hd__a22o_1 _15415_ (.A1(_10365_),
    .A2(\line_cache[108][3] ),
    .B1(_10366_),
    .B2(\line_cache[109][3] ),
    .X(_11138_));
 sky130_fd_sc_hd__a221o_1 _15416_ (.A1(\line_cache[111][3] ),
    .A2(_10363_),
    .B1(\line_cache[110][3] ),
    .B2(_10364_),
    .C1(_11138_),
    .X(_11139_));
 sky130_fd_sc_hd__or2_1 _15417_ (.A(_11137_),
    .B(_11139_),
    .X(_11140_));
 sky130_fd_sc_hd__or4_1 _15418_ (.A(_11129_),
    .B(_11130_),
    .C(_11132_),
    .D(_11140_),
    .X(_11141_));
 sky130_fd_sc_hd__nor2_1 _15419_ (.A(_11128_),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__and3_1 _15420_ (.A(_10176_),
    .B(\line_cache[121][3] ),
    .C(_10302_),
    .X(_11143_));
 sky130_fd_sc_hd__a21o_1 _15421_ (.A1(\line_cache[120][3] ),
    .A2(_10317_),
    .B1(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__a221o_1 _15422_ (.A1(\line_cache[123][3] ),
    .A2(_10315_),
    .B1(\line_cache[122][3] ),
    .B2(_10316_),
    .C1(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__a22o_1 _15423_ (.A1(_10298_),
    .A2(\line_cache[112][3] ),
    .B1(_10299_),
    .B2(\line_cache[113][3] ),
    .X(_11146_));
 sky130_fd_sc_hd__a221o_1 _15424_ (.A1(\line_cache[115][3] ),
    .A2(_10296_),
    .B1(\line_cache[114][3] ),
    .B2(_10297_),
    .C1(_11146_),
    .X(_11147_));
 sky130_fd_sc_hd__a22o_1 _15425_ (.A1(_10311_),
    .A2(\line_cache[116][3] ),
    .B1(_10312_),
    .B2(\line_cache[117][3] ),
    .X(_11148_));
 sky130_fd_sc_hd__a221o_1 _15426_ (.A1(\line_cache[119][3] ),
    .A2(_10309_),
    .B1(\line_cache[118][3] ),
    .B2(_10310_),
    .C1(_11148_),
    .X(_11149_));
 sky130_fd_sc_hd__a22o_1 _15427_ (.A1(_10305_),
    .A2(\line_cache[124][3] ),
    .B1(_10306_),
    .B2(\line_cache[125][3] ),
    .X(_11150_));
 sky130_fd_sc_hd__a221o_1 _15428_ (.A1(\line_cache[126][3] ),
    .A2(_10304_),
    .B1(\line_cache[127][3] ),
    .B2(_10622_),
    .C1(_11150_),
    .X(_11151_));
 sky130_fd_sc_hd__or4_1 _15429_ (.A(_11145_),
    .B(_11147_),
    .C(_11149_),
    .D(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__and3_1 _15430_ (.A(_09758_),
    .B(_10098_),
    .C(\line_cache[133][3] ),
    .X(_11153_));
 sky130_fd_sc_hd__a21o_1 _15431_ (.A1(\line_cache[132][3] ),
    .A2(_10324_),
    .B1(_11153_),
    .X(_11154_));
 sky130_fd_sc_hd__a221o_1 _15432_ (.A1(\line_cache[135][3] ),
    .A2(_10322_),
    .B1(\line_cache[134][3] ),
    .B2(_10323_),
    .C1(_11154_),
    .X(_11155_));
 sky130_fd_sc_hd__and3_1 _15433_ (.A(_09758_),
    .B(_10031_),
    .C(\line_cache[141][3] ),
    .X(_11156_));
 sky130_fd_sc_hd__a21o_1 _15434_ (.A1(\line_cache[140][3] ),
    .A2(_10336_),
    .B1(_11156_),
    .X(_11157_));
 sky130_fd_sc_hd__a221o_1 _15435_ (.A1(\line_cache[143][3] ),
    .A2(_10334_),
    .B1(\line_cache[142][3] ),
    .B2(_10335_),
    .C1(_11157_),
    .X(_11158_));
 sky130_fd_sc_hd__a22o_1 _15436_ (.A1(_10330_),
    .A2(\line_cache[129][3] ),
    .B1(\line_cache[128][3] ),
    .B2(_10629_),
    .X(_11159_));
 sky130_fd_sc_hd__a221o_1 _15437_ (.A1(\line_cache[131][3] ),
    .A2(_10328_),
    .B1(\line_cache[130][3] ),
    .B2(_10329_),
    .C1(_11159_),
    .X(_11160_));
 sky130_fd_sc_hd__a22o_1 _15438_ (.A1(_10342_),
    .A2(\line_cache[139][3] ),
    .B1(\line_cache[138][3] ),
    .B2(_10343_),
    .X(_11161_));
 sky130_fd_sc_hd__a221o_1 _15439_ (.A1(\line_cache[137][3] ),
    .A2(_10340_),
    .B1(\line_cache[136][3] ),
    .B2(_10341_),
    .C1(_11161_),
    .X(_11162_));
 sky130_fd_sc_hd__or4_2 _15440_ (.A(_11155_),
    .B(_11158_),
    .C(_11160_),
    .D(_11162_),
    .X(_11163_));
 sky130_fd_sc_hd__nor2_1 _15441_ (.A(_11152_),
    .B(_11163_),
    .Y(_11164_));
 sky130_fd_sc_hd__and3_2 _15442_ (.A(_11119_),
    .B(_11142_),
    .C(_11164_),
    .X(_11165_));
 sky130_fd_sc_hd__nand3_1 _15443_ (.A(_11024_),
    .B(_11087_),
    .C(_11165_),
    .Y(_11166_));
 sky130_fd_sc_hd__o21ba_2 _15444_ (.A1(_10915_),
    .A2(_11166_),
    .B1_N(_08979_),
    .X(_11167_));
 sky130_fd_sc_hd__buf_6 _15445_ (.A(_11167_),
    .X(net129));
 sky130_fd_sc_hd__and2_1 _15446_ (.A(_09912_),
    .B(\line_cache[0][4] ),
    .X(_11168_));
 sky130_fd_sc_hd__and3_1 _15447_ (.A(_10031_),
    .B(\line_cache[77][4] ),
    .C(_10167_),
    .X(_11169_));
 sky130_fd_sc_hd__and3_1 _15448_ (.A(_10038_),
    .B(\line_cache[78][4] ),
    .C(_10167_),
    .X(_11170_));
 sky130_fd_sc_hd__and3_1 _15449_ (.A(_10041_),
    .B(\line_cache[76][4] ),
    .C(_10161_),
    .X(_11171_));
 sky130_fd_sc_hd__a2111o_1 _15450_ (.A1(_10168_),
    .A2(\line_cache[79][4] ),
    .B1(_11169_),
    .C1(_11170_),
    .D1(_11171_),
    .X(_11172_));
 sky130_fd_sc_hd__a22o_1 _15451_ (.A1(_10182_),
    .A2(\line_cache[64][4] ),
    .B1(_10183_),
    .B2(\line_cache[65][4] ),
    .X(_11173_));
 sky130_fd_sc_hd__a221o_1 _15452_ (.A1(\line_cache[67][4] ),
    .A2(_10180_),
    .B1(\line_cache[66][4] ),
    .B2(_10181_),
    .C1(_11173_),
    .X(_11174_));
 sky130_fd_sc_hd__a22o_1 _15453_ (.A1(_10163_),
    .A2(\line_cache[68][4] ),
    .B1(_10164_),
    .B2(\line_cache[69][4] ),
    .X(_11175_));
 sky130_fd_sc_hd__a221o_1 _15454_ (.A1(\line_cache[71][4] ),
    .A2(_10159_),
    .B1(\line_cache[70][4] ),
    .B2(_10750_),
    .C1(_11175_),
    .X(_11176_));
 sky130_fd_sc_hd__a22o_1 _15455_ (.A1(_10175_),
    .A2(\line_cache[72][4] ),
    .B1(_10753_),
    .B2(\line_cache[73][4] ),
    .X(_11177_));
 sky130_fd_sc_hd__a221o_1 _15456_ (.A1(\line_cache[75][4] ),
    .A2(_10173_),
    .B1(\line_cache[74][4] ),
    .B2(_10174_),
    .C1(_11177_),
    .X(_11178_));
 sky130_fd_sc_hd__or4_4 _15457_ (.A(_11172_),
    .B(_11174_),
    .C(_11176_),
    .D(_11178_),
    .X(_11179_));
 sky130_fd_sc_hd__a22o_1 _15458_ (.A1(_10189_),
    .A2(\line_cache[252][4] ),
    .B1(_10190_),
    .B2(\line_cache[251][4] ),
    .X(_11180_));
 sky130_fd_sc_hd__a221o_1 _15459_ (.A1(\line_cache[254][4] ),
    .A2(_10187_),
    .B1(\line_cache[253][4] ),
    .B2(_10188_),
    .C1(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__a22o_1 _15460_ (.A1(_10195_),
    .A2(\line_cache[248][4] ),
    .B1(_10196_),
    .B2(\line_cache[247][4] ),
    .X(_11182_));
 sky130_fd_sc_hd__a221o_1 _15461_ (.A1(\line_cache[250][4] ),
    .A2(_10193_),
    .B1(\line_cache[249][4] ),
    .B2(_10194_),
    .C1(_11182_),
    .X(_11183_));
 sky130_fd_sc_hd__and2b_1 _15462_ (.A_N(_10200_),
    .B(\line_cache[240][4] ),
    .X(_11184_));
 sky130_fd_sc_hd__and2b_1 _15463_ (.A_N(_09570_),
    .B(\line_cache[241][4] ),
    .X(_11185_));
 sky130_fd_sc_hd__and2b_1 _15464_ (.A_N(_10203_),
    .B(\line_cache[242][4] ),
    .X(_11186_));
 sky130_fd_sc_hd__a2111o_1 _15465_ (.A1(\line_cache[239][4] ),
    .A2(_10199_),
    .B1(_11184_),
    .C1(_11185_),
    .D1(_11186_),
    .X(_11187_));
 sky130_fd_sc_hd__and2b_1 _15466_ (.A_N(_10206_),
    .B(\line_cache[243][4] ),
    .X(_11188_));
 sky130_fd_sc_hd__and2b_1 _15467_ (.A_N(_10208_),
    .B(\line_cache[244][4] ),
    .X(_11189_));
 sky130_fd_sc_hd__and2b_1 _15468_ (.A_N(_09597_),
    .B(\line_cache[245][4] ),
    .X(_11190_));
 sky130_fd_sc_hd__and2b_1 _15469_ (.A_N(_10211_),
    .B(\line_cache[246][4] ),
    .X(_11191_));
 sky130_fd_sc_hd__or4_1 _15470_ (.A(_11188_),
    .B(_11189_),
    .C(_11190_),
    .D(_11191_),
    .X(_11192_));
 sky130_fd_sc_hd__or4_1 _15471_ (.A(_11181_),
    .B(_11183_),
    .C(_11187_),
    .D(_11192_),
    .X(_11193_));
 sky130_fd_sc_hd__and3_1 _15472_ (.A(_09595_),
    .B(\line_cache[229][4] ),
    .C(_10099_),
    .X(_11194_));
 sky130_fd_sc_hd__and3_1 _15473_ (.A(_10044_),
    .B(\line_cache[230][4] ),
    .C(_10434_),
    .X(_11195_));
 sky130_fd_sc_hd__and3_1 _15474_ (.A(_10104_),
    .B(\line_cache[227][4] ),
    .C(_10434_),
    .X(_11196_));
 sky130_fd_sc_hd__and3_1 _15475_ (.A(_10106_),
    .B(\line_cache[228][4] ),
    .C(_10437_),
    .X(_11197_));
 sky130_fd_sc_hd__or4_1 _15476_ (.A(_11194_),
    .B(_11195_),
    .C(_11196_),
    .D(_11197_),
    .X(_11198_));
 sky130_fd_sc_hd__and3_1 _15477_ (.A(_09544_),
    .B(\line_cache[223][4] ),
    .C(_10109_),
    .X(_11199_));
 sky130_fd_sc_hd__and3_1 _15478_ (.A(_10070_),
    .B(\line_cache[224][4] ),
    .C(_10434_),
    .X(_11200_));
 sky130_fd_sc_hd__and3_1 _15479_ (.A(_10067_),
    .B(\line_cache[225][4] ),
    .C(_10437_),
    .X(_11201_));
 sky130_fd_sc_hd__and3_1 _15480_ (.A(_10074_),
    .B(\line_cache[226][4] ),
    .C(_10437_),
    .X(_11202_));
 sky130_fd_sc_hd__or4_1 _15481_ (.A(_11199_),
    .B(_11200_),
    .C(_11201_),
    .D(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__a22o_1 _15482_ (.A1(_10118_),
    .A2(\line_cache[236][4] ),
    .B1(_10120_),
    .B2(\line_cache[235][4] ),
    .X(_11204_));
 sky130_fd_sc_hd__a221o_1 _15483_ (.A1(\line_cache[238][4] ),
    .A2(_10116_),
    .B1(\line_cache[237][4] ),
    .B2(_10117_),
    .C1(_11204_),
    .X(_11205_));
 sky130_fd_sc_hd__a22o_1 _15484_ (.A1(_10125_),
    .A2(\line_cache[232][4] ),
    .B1(_10126_),
    .B2(\line_cache[231][4] ),
    .X(_11206_));
 sky130_fd_sc_hd__a221o_1 _15485_ (.A1(\line_cache[234][4] ),
    .A2(_10123_),
    .B1(\line_cache[233][4] ),
    .B2(_10124_),
    .C1(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__or4_1 _15486_ (.A(_11198_),
    .B(_11203_),
    .C(_11205_),
    .D(_11207_),
    .X(_11208_));
 sky130_fd_sc_hd__a22o_1 _15487_ (.A1(_10132_),
    .A2(\line_cache[220][4] ),
    .B1(_10133_),
    .B2(\line_cache[219][4] ),
    .X(_11209_));
 sky130_fd_sc_hd__a221o_1 _15488_ (.A1(\line_cache[222][4] ),
    .A2(_10130_),
    .B1(\line_cache[221][4] ),
    .B2(_10131_),
    .C1(_11209_),
    .X(_11210_));
 sky130_fd_sc_hd__a22o_1 _15489_ (.A1(_10138_),
    .A2(\line_cache[208][4] ),
    .B1(_10139_),
    .B2(\line_cache[207][4] ),
    .X(_11211_));
 sky130_fd_sc_hd__a221o_1 _15490_ (.A1(\line_cache[210][4] ),
    .A2(_10136_),
    .B1(\line_cache[209][4] ),
    .B2(_10137_),
    .C1(_11211_),
    .X(_11212_));
 sky130_fd_sc_hd__a22o_1 _15491_ (.A1(_10144_),
    .A2(\line_cache[216][4] ),
    .B1(_10145_),
    .B2(\line_cache[215][4] ),
    .X(_11213_));
 sky130_fd_sc_hd__a221o_1 _15492_ (.A1(\line_cache[218][4] ),
    .A2(_10142_),
    .B1(\line_cache[217][4] ),
    .B2(_10143_),
    .C1(_11213_),
    .X(_11214_));
 sky130_fd_sc_hd__and2b_1 _15493_ (.A_N(_10148_),
    .B(\line_cache[211][4] ),
    .X(_11215_));
 sky130_fd_sc_hd__nor2b_1 _15494_ (.A(_10150_),
    .B_N(\line_cache[212][4] ),
    .Y(_11216_));
 sky130_fd_sc_hd__and2b_1 _15495_ (.A_N(_10152_),
    .B(\line_cache[213][4] ),
    .X(_11217_));
 sky130_fd_sc_hd__and2b_1 _15496_ (.A_N(_10154_),
    .B(\line_cache[214][4] ),
    .X(_11218_));
 sky130_fd_sc_hd__or4_1 _15497_ (.A(_11215_),
    .B(_11216_),
    .C(_11217_),
    .D(_11218_),
    .X(_11219_));
 sky130_fd_sc_hd__or4_2 _15498_ (.A(_11210_),
    .B(_11212_),
    .C(_11214_),
    .D(_11219_),
    .X(_11220_));
 sky130_fd_sc_hd__or2_1 _15499_ (.A(_11208_),
    .B(_11220_),
    .X(_11221_));
 sky130_fd_sc_hd__or3_1 _15500_ (.A(_11179_),
    .B(_11193_),
    .C(_11221_),
    .X(_11222_));
 sky130_fd_sc_hd__and3_1 _15501_ (.A(_10035_),
    .B(\line_cache[203][4] ),
    .C(_09539_),
    .X(_11223_));
 sky130_fd_sc_hd__and3_1 _15502_ (.A(_10038_),
    .B(\line_cache[206][4] ),
    .C(_10075_),
    .X(_11224_));
 sky130_fd_sc_hd__and3_1 _15503_ (.A(_10041_),
    .B(\line_cache[204][4] ),
    .C(_10075_),
    .X(_11225_));
 sky130_fd_sc_hd__a2111o_1 _15504_ (.A1(\line_cache[205][4] ),
    .A2(_10033_),
    .B1(_11223_),
    .C1(_11224_),
    .D1(_11225_),
    .X(_11226_));
 sky130_fd_sc_hd__a22o_1 _15505_ (.A1(_10049_),
    .A2(\line_cache[195][4] ),
    .B1(\line_cache[196][4] ),
    .B2(_10051_),
    .X(_11227_));
 sky130_fd_sc_hd__a221o_1 _15506_ (.A1(\line_cache[198][4] ),
    .A2(_10046_),
    .B1(\line_cache[197][4] ),
    .B2(_10047_),
    .C1(_11227_),
    .X(_11228_));
 sky130_fd_sc_hd__a22o_1 _15507_ (.A1(_10060_),
    .A2(\line_cache[200][4] ),
    .B1(_10063_),
    .B2(\line_cache[199][4] ),
    .X(_11229_));
 sky130_fd_sc_hd__a221o_1 _15508_ (.A1(\line_cache[202][4] ),
    .A2(_10056_),
    .B1(\line_cache[201][4] ),
    .B2(_10059_),
    .C1(_11229_),
    .X(_11230_));
 sky130_fd_sc_hd__and3_1 _15509_ (.A(_10067_),
    .B(\line_cache[193][4] ),
    .C(_09540_),
    .X(_11231_));
 sky130_fd_sc_hd__and3_1 _15510_ (.A(_10071_),
    .B(\line_cache[192][4] ),
    .C(_09540_),
    .X(_11232_));
 sky130_fd_sc_hd__and3_1 _15511_ (.A(_10074_),
    .B(\line_cache[194][4] ),
    .C(_09540_),
    .X(_11233_));
 sky130_fd_sc_hd__a2111o_1 _15512_ (.A1(_10066_),
    .A2(\line_cache[286][4] ),
    .B1(_11231_),
    .C1(_11232_),
    .D1(_11233_),
    .X(_11234_));
 sky130_fd_sc_hd__or4_1 _15513_ (.A(_11226_),
    .B(_11228_),
    .C(_11230_),
    .D(_11234_),
    .X(_11235_));
 sky130_fd_sc_hd__a22o_1 _15514_ (.A1(_09623_),
    .A2(\line_cache[275][4] ),
    .B1(_09620_),
    .B2(\line_cache[274][4] ),
    .X(_11236_));
 sky130_fd_sc_hd__a22o_1 _15515_ (.A1(_10080_),
    .A2(\line_cache[276][4] ),
    .B1(\line_cache[277][4] ),
    .B2(_10081_),
    .X(_11237_));
 sky130_fd_sc_hd__a22o_1 _15516_ (.A1(_10086_),
    .A2(\line_cache[270][4] ),
    .B1(\line_cache[269][4] ),
    .B2(_10088_),
    .X(_11238_));
 sky130_fd_sc_hd__a221o_1 _15517_ (.A1(\line_cache[273][4] ),
    .A2(_10083_),
    .B1(\line_cache[272][4] ),
    .B2(_10084_),
    .C1(_11238_),
    .X(_11239_));
 sky130_fd_sc_hd__a22o_1 _15518_ (.A1(_09658_),
    .A2(\line_cache[283][4] ),
    .B1(\line_cache[282][4] ),
    .B2(_09661_),
    .X(_11240_));
 sky130_fd_sc_hd__a22o_1 _15519_ (.A1(_09645_),
    .A2(\line_cache[285][4] ),
    .B1(\line_cache[284][4] ),
    .B2(_09648_),
    .X(_11241_));
 sky130_fd_sc_hd__a22o_1 _15520_ (.A1(_09639_),
    .A2(\line_cache[279][4] ),
    .B1(\line_cache[278][4] ),
    .B2(_09636_),
    .X(_11242_));
 sky130_fd_sc_hd__a221o_1 _15521_ (.A1(\line_cache[281][4] ),
    .A2(_09663_),
    .B1(\line_cache[280][4] ),
    .B2(_09655_),
    .C1(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__or3_1 _15522_ (.A(_11240_),
    .B(_11241_),
    .C(_11243_),
    .X(_11244_));
 sky130_fd_sc_hd__or4_1 _15523_ (.A(_11236_),
    .B(_11237_),
    .C(_11239_),
    .D(_11244_),
    .X(_11245_));
 sky130_fd_sc_hd__nor2_1 _15524_ (.A(_11235_),
    .B(_11245_),
    .Y(_11246_));
 sky130_fd_sc_hd__and2b_1 _15525_ (.A_N(_09987_),
    .B(\line_cache[256][4] ),
    .X(_11247_));
 sky130_fd_sc_hd__and2b_1 _15526_ (.A_N(_09747_),
    .B(\line_cache[302][4] ),
    .X(_11248_));
 sky130_fd_sc_hd__a22o_1 _15527_ (.A1(_09743_),
    .A2(\line_cache[301][4] ),
    .B1(\line_cache[300][4] ),
    .B2(_09742_),
    .X(_11249_));
 sky130_fd_sc_hd__or3_1 _15528_ (.A(_11247_),
    .B(_11248_),
    .C(_11249_),
    .X(_11250_));
 sky130_fd_sc_hd__and3_1 _15529_ (.A(_09917_),
    .B(_09691_),
    .C(\line_cache[258][4] ),
    .X(_11251_));
 sky130_fd_sc_hd__and3_1 _15530_ (.A(_09848_),
    .B(_09691_),
    .C(\line_cache[260][4] ),
    .X(_11252_));
 sky130_fd_sc_hd__and3_1 _15531_ (.A(_09919_),
    .B(_09611_),
    .C(\line_cache[257][4] ),
    .X(_11253_));
 sky130_fd_sc_hd__and3_1 _15532_ (.A(_09840_),
    .B(_09611_),
    .C(\line_cache[259][4] ),
    .X(_11254_));
 sky130_fd_sc_hd__or4_1 _15533_ (.A(_11251_),
    .B(_11252_),
    .C(_11253_),
    .D(_11254_),
    .X(_11255_));
 sky130_fd_sc_hd__and3_1 _15534_ (.A(_09858_),
    .B(_09547_),
    .C(\line_cache[267][4] ),
    .X(_11256_));
 sky130_fd_sc_hd__a22o_1 _15535_ (.A1(_09998_),
    .A2(\line_cache[265][4] ),
    .B1(\line_cache[266][4] ),
    .B2(_09999_),
    .X(_11257_));
 sky130_fd_sc_hd__a311o_1 _15536_ (.A1(_09548_),
    .A2(\line_cache[268][4] ),
    .A3(_09862_),
    .B1(_11256_),
    .C1(_11257_),
    .X(_11258_));
 sky130_fd_sc_hd__nand2_1 _15537_ (.A(_10007_),
    .B(\line_cache[262][4] ),
    .Y(_11259_));
 sky130_fd_sc_hd__nand2_1 _15538_ (.A(_10010_),
    .B(\line_cache[261][4] ),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_1 _15539_ (.A(_11259_),
    .B(_11260_),
    .Y(_11261_));
 sky130_fd_sc_hd__a221oi_1 _15540_ (.A1(_10003_),
    .A2(\line_cache[264][4] ),
    .B1(_10005_),
    .B2(\line_cache[263][4] ),
    .C1(_11261_),
    .Y(_11262_));
 sky130_fd_sc_hd__or4b_1 _15541_ (.A(_11250_),
    .B(_11255_),
    .C(_11258_),
    .D_N(_11262_),
    .X(_11263_));
 sky130_fd_sc_hd__a22o_1 _15542_ (.A1(_09682_),
    .A2(\line_cache[308][4] ),
    .B1(\line_cache[309][4] ),
    .B2(_09685_),
    .X(_11264_));
 sky130_fd_sc_hd__a221o_1 _15543_ (.A1(\line_cache[311][4] ),
    .A2(_09689_),
    .B1(\line_cache[310][4] ),
    .B2(_09693_),
    .C1(_11264_),
    .X(_11265_));
 sky130_fd_sc_hd__a22o_1 _15544_ (.A1(_09728_),
    .A2(\line_cache[295][4] ),
    .B1(\line_cache[294][4] ),
    .B2(_09726_),
    .X(_11266_));
 sky130_fd_sc_hd__a221o_1 _15545_ (.A1(\line_cache[293][4] ),
    .A2(_09730_),
    .B1(\line_cache[292][4] ),
    .B2(_10018_),
    .C1(_11266_),
    .X(_11267_));
 sky130_fd_sc_hd__a22o_1 _15546_ (.A1(_09716_),
    .A2(\line_cache[296][4] ),
    .B1(\line_cache[297][4] ),
    .B2(_09721_),
    .X(_11268_));
 sky130_fd_sc_hd__a221o_1 _15547_ (.A1(\line_cache[299][4] ),
    .A2(_09718_),
    .B1(\line_cache[298][4] ),
    .B2(_09720_),
    .C1(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__a22o_1 _15548_ (.A1(_10025_),
    .A2(\line_cache[288][4] ),
    .B1(\line_cache[289][4] ),
    .B2(_10026_),
    .X(_11270_));
 sky130_fd_sc_hd__a221o_1 _15549_ (.A1(\line_cache[291][4] ),
    .A2(_10023_),
    .B1(\line_cache[290][4] ),
    .B2(_10024_),
    .C1(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__or4_4 _15550_ (.A(_11265_),
    .B(_11267_),
    .C(_11269_),
    .D(_11271_),
    .X(_11272_));
 sky130_fd_sc_hd__nor2_1 _15551_ (.A(_11263_),
    .B(_11272_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand2_1 _15552_ (.A(_11246_),
    .B(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_11222_),
    .B(_11274_),
    .Y(_11275_));
 sky130_fd_sc_hd__a22o_1 _15554_ (.A1(_09842_),
    .A2(\line_cache[6][4] ),
    .B1(\line_cache[5][4] ),
    .B2(_09844_),
    .X(_11276_));
 sky130_fd_sc_hd__a221o_1 _15555_ (.A1(\line_cache[4][4] ),
    .A2(_09850_),
    .B1(\line_cache[3][4] ),
    .B2(_09914_),
    .C1(_11276_),
    .X(_11277_));
 sky130_fd_sc_hd__and3_1 _15556_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][4] ),
    .X(_11278_));
 sky130_fd_sc_hd__and3_1 _15557_ (.A(_09919_),
    .B(_09533_),
    .C(\line_cache[1][4] ),
    .X(_11279_));
 sky130_fd_sc_hd__a211o_1 _15558_ (.A1(\line_cache[15][4] ),
    .A2(_09867_),
    .B1(_11278_),
    .C1(_11279_),
    .X(_11280_));
 sky130_fd_sc_hd__and3_1 _15559_ (.A(_09922_),
    .B(_09532_),
    .C(\line_cache[63][4] ),
    .X(_11281_));
 sky130_fd_sc_hd__a31o_1 _15560_ (.A1(_09548_),
    .A2(\line_cache[319][4] ),
    .A3(_09922_),
    .B1(_11281_),
    .X(_11282_));
 sky130_fd_sc_hd__a221o_1 _15561_ (.A1(\line_cache[47][4] ),
    .A2(_09806_),
    .B1(\line_cache[31][4] ),
    .B2(_09907_),
    .C1(_11282_),
    .X(_11283_));
 sky130_fd_sc_hd__nand2_1 _15562_ (.A(_09746_),
    .B(\line_cache[303][4] ),
    .Y(_11284_));
 sky130_fd_sc_hd__nand2_1 _15563_ (.A(_09930_),
    .B(\line_cache[271][4] ),
    .Y(_11285_));
 sky130_fd_sc_hd__nand2_1 _15564_ (.A(_11284_),
    .B(_11285_),
    .Y(_11286_));
 sky130_fd_sc_hd__a221oi_2 _15565_ (.A1(\line_cache[255][4] ),
    .A2(_09926_),
    .B1(\line_cache[287][4] ),
    .B2(_09927_),
    .C1(_11286_),
    .Y(_11287_));
 sky130_fd_sc_hd__or4b_1 _15566_ (.A(_11277_),
    .B(_11280_),
    .C(_11283_),
    .D_N(_11287_),
    .X(_11288_));
 sky130_fd_sc_hd__a22o_1 _15567_ (.A1(_09803_),
    .A2(\line_cache[45][4] ),
    .B1(\line_cache[46][4] ),
    .B2(_09804_),
    .X(_11289_));
 sky130_fd_sc_hd__a22o_1 _15568_ (.A1(_09824_),
    .A2(\line_cache[48][4] ),
    .B1(\line_cache[49][4] ),
    .B2(_09826_),
    .X(_11290_));
 sky130_fd_sc_hd__nand2_1 _15569_ (.A(_09787_),
    .B(\line_cache[41][4] ),
    .Y(_11291_));
 sky130_fd_sc_hd__nand2_1 _15570_ (.A(_09789_),
    .B(\line_cache[42][4] ),
    .Y(_11292_));
 sky130_fd_sc_hd__nand2_1 _15571_ (.A(_11291_),
    .B(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__a221oi_2 _15572_ (.A1(_09785_),
    .A2(\line_cache[43][4] ),
    .B1(\line_cache[44][4] ),
    .B2(_09801_),
    .C1(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__or3b_1 _15573_ (.A(_11289_),
    .B(_11290_),
    .C_N(_11294_),
    .X(_11295_));
 sky130_fd_sc_hd__a22o_1 _15574_ (.A1(_09699_),
    .A2(\line_cache[317][4] ),
    .B1(\line_cache[316][4] ),
    .B2(_09697_),
    .X(_11296_));
 sky130_fd_sc_hd__a22o_1 _15575_ (.A1(_09832_),
    .A2(\line_cache[58][4] ),
    .B1(\line_cache[59][4] ),
    .B2(_09833_),
    .X(_11297_));
 sky130_fd_sc_hd__a22o_1 _15576_ (.A1(_09819_),
    .A2(\line_cache[61][4] ),
    .B1(\line_cache[60][4] ),
    .B2(_09817_),
    .X(_11298_));
 sky130_fd_sc_hd__a22o_1 _15577_ (.A1(_09822_),
    .A2(\line_cache[62][4] ),
    .B1(\line_cache[318][4] ),
    .B2(_09702_),
    .X(_11299_));
 sky130_fd_sc_hd__or4_1 _15578_ (.A(_11296_),
    .B(_11297_),
    .C(_11298_),
    .D(_11299_),
    .X(_11300_));
 sky130_fd_sc_hd__a22o_1 _15579_ (.A1(_09675_),
    .A2(\line_cache[304][4] ),
    .B1(\line_cache[305][4] ),
    .B2(_09676_),
    .X(_11301_));
 sky130_fd_sc_hd__a22o_1 _15580_ (.A1(_09705_),
    .A2(\line_cache[312][4] ),
    .B1(\line_cache[313][4] ),
    .B2(_09707_),
    .X(_11302_));
 sky130_fd_sc_hd__a22o_1 _15581_ (.A1(_09708_),
    .A2(\line_cache[314][4] ),
    .B1(\line_cache[315][4] ),
    .B2(_09709_),
    .X(_11303_));
 sky130_fd_sc_hd__a22o_1 _15582_ (.A1(_09677_),
    .A2(\line_cache[306][4] ),
    .B1(\line_cache[307][4] ),
    .B2(_09678_),
    .X(_11304_));
 sky130_fd_sc_hd__or4_1 _15583_ (.A(_11301_),
    .B(_11302_),
    .C(_11303_),
    .D(_11304_),
    .X(_11305_));
 sky130_fd_sc_hd__a22o_1 _15584_ (.A1(_09830_),
    .A2(\line_cache[56][4] ),
    .B1(\line_cache[57][4] ),
    .B2(_09834_),
    .X(_11306_));
 sky130_fd_sc_hd__a22o_1 _15585_ (.A1(_09809_),
    .A2(\line_cache[52][4] ),
    .B1(\line_cache[53][4] ),
    .B2(_09811_),
    .X(_11307_));
 sky130_fd_sc_hd__a22o_1 _15586_ (.A1(_09827_),
    .A2(\line_cache[50][4] ),
    .B1(\line_cache[51][4] ),
    .B2(_09828_),
    .X(_11308_));
 sky130_fd_sc_hd__a22o_1 _15587_ (.A1(_09813_),
    .A2(\line_cache[54][4] ),
    .B1(\line_cache[55][4] ),
    .B2(_09815_),
    .X(_11309_));
 sky130_fd_sc_hd__or4_1 _15588_ (.A(_11306_),
    .B(_11307_),
    .C(_11308_),
    .D(_11309_),
    .X(_11310_));
 sky130_fd_sc_hd__or4_2 _15589_ (.A(_11295_),
    .B(_11300_),
    .C(_11305_),
    .D(_11310_),
    .X(_11311_));
 sky130_fd_sc_hd__nand2_1 _15590_ (.A(_09864_),
    .B(\line_cache[12][4] ),
    .Y(_11312_));
 sky130_fd_sc_hd__nand2_1 _15591_ (.A(_09860_),
    .B(\line_cache[11][4] ),
    .Y(_11313_));
 sky130_fd_sc_hd__nand2_1 _15592_ (.A(_11312_),
    .B(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__a221oi_2 _15593_ (.A1(_09870_),
    .A2(\line_cache[14][4] ),
    .B1(\line_cache[13][4] ),
    .B2(_09873_),
    .C1(_11314_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_1 _15594_ (.A(_09853_),
    .B(\line_cache[10][4] ),
    .Y(_11316_));
 sky130_fd_sc_hd__nand2_1 _15595_ (.A(_09857_),
    .B(\line_cache[9][4] ),
    .Y(_11317_));
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(_11316_),
    .B(_11317_),
    .Y(_11318_));
 sky130_fd_sc_hd__a221oi_1 _15597_ (.A1(_09855_),
    .A2(\line_cache[8][4] ),
    .B1(_09847_),
    .B2(\line_cache[7][4] ),
    .C1(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__nand2_1 _15598_ (.A(_11315_),
    .B(_11319_),
    .Y(_11320_));
 sky130_fd_sc_hd__and3_1 _15599_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][4] ),
    .X(_11321_));
 sky130_fd_sc_hd__a22o_1 _15600_ (.A1(_09884_),
    .A2(\line_cache[23][4] ),
    .B1(\line_cache[22][4] ),
    .B2(_09886_),
    .X(_11322_));
 sky130_fd_sc_hd__a22o_1 _15601_ (.A1(_09877_),
    .A2(\line_cache[19][4] ),
    .B1(\line_cache[18][4] ),
    .B2(_09878_),
    .X(_11323_));
 sky130_fd_sc_hd__a221o_1 _15602_ (.A1(\line_cache[17][4] ),
    .A2(_09969_),
    .B1(\line_cache[16][4] ),
    .B2(_09970_),
    .C1(_11323_),
    .X(_11324_));
 sky130_fd_sc_hd__a2111o_1 _15603_ (.A1(\line_cache[20][4] ),
    .A2(_09888_),
    .B1(_11321_),
    .C1(_11322_),
    .D1(_11324_),
    .X(_11325_));
 sky130_fd_sc_hd__a22o_1 _15604_ (.A1(_09796_),
    .A2(\line_cache[33][4] ),
    .B1(\line_cache[34][4] ),
    .B2(_09798_),
    .X(_11326_));
 sky130_fd_sc_hd__a221o_1 _15605_ (.A1(\line_cache[36][4] ),
    .A2(_09777_),
    .B1(\line_cache[35][4] ),
    .B2(_09794_),
    .C1(_11326_),
    .X(_11327_));
 sky130_fd_sc_hd__a22o_1 _15606_ (.A1(_09890_),
    .A2(\line_cache[27][4] ),
    .B1(\line_cache[26][4] ),
    .B2(_09896_),
    .X(_11328_));
 sky130_fd_sc_hd__a221oi_2 _15607_ (.A1(\line_cache[25][4] ),
    .A2(_09892_),
    .B1(\line_cache[24][4] ),
    .B2(_09895_),
    .C1(_11328_),
    .Y(_11329_));
 sky130_fd_sc_hd__a22o_1 _15608_ (.A1(_09903_),
    .A2(\line_cache[29][4] ),
    .B1(\line_cache[28][4] ),
    .B2(_09900_),
    .X(_11330_));
 sky130_fd_sc_hd__a221oi_1 _15609_ (.A1(\line_cache[32][4] ),
    .A2(_09792_),
    .B1(\line_cache[30][4] ),
    .B2(_09905_),
    .C1(_11330_),
    .Y(_11331_));
 sky130_fd_sc_hd__nand2_1 _15610_ (.A(_09773_),
    .B(\line_cache[38][4] ),
    .Y(_11332_));
 sky130_fd_sc_hd__nand2_1 _15611_ (.A(_09775_),
    .B(\line_cache[37][4] ),
    .Y(_11333_));
 sky130_fd_sc_hd__nand2_1 _15612_ (.A(_11332_),
    .B(_11333_),
    .Y(_11334_));
 sky130_fd_sc_hd__a221oi_2 _15613_ (.A1(_09783_),
    .A2(\line_cache[40][4] ),
    .B1(\line_cache[39][4] ),
    .B2(_09780_),
    .C1(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__and4b_1 _15614_ (.A_N(_11327_),
    .B(_11329_),
    .C(_11331_),
    .D(_11335_),
    .X(_11336_));
 sky130_fd_sc_hd__or3b_2 _15615_ (.A(_11320_),
    .B(_11325_),
    .C_N(_11336_),
    .X(_11337_));
 sky130_fd_sc_hd__nor3_2 _15616_ (.A(_11288_),
    .B(_11311_),
    .C(_11337_),
    .Y(_11338_));
 sky130_fd_sc_hd__a22o_1 _15617_ (.A1(_10378_),
    .A2(\line_cache[80][4] ),
    .B1(_10379_),
    .B2(\line_cache[81][4] ),
    .X(_11339_));
 sky130_fd_sc_hd__a221o_1 _15618_ (.A1(\line_cache[83][4] ),
    .A2(_10376_),
    .B1(\line_cache[82][4] ),
    .B2(_10377_),
    .C1(_11339_),
    .X(_11340_));
 sky130_fd_sc_hd__a22o_1 _15619_ (.A1(_10384_),
    .A2(\line_cache[92][4] ),
    .B1(_10385_),
    .B2(\line_cache[93][4] ),
    .X(_11341_));
 sky130_fd_sc_hd__a221o_1 _15620_ (.A1(\line_cache[95][4] ),
    .A2(net136),
    .B1(\line_cache[94][4] ),
    .B2(_10383_),
    .C1(_11341_),
    .X(_11342_));
 sky130_fd_sc_hd__a22o_1 _15621_ (.A1(_10390_),
    .A2(\line_cache[84][4] ),
    .B1(_10391_),
    .B2(\line_cache[85][4] ),
    .X(_11343_));
 sky130_fd_sc_hd__a221o_1 _15622_ (.A1(\line_cache[87][4] ),
    .A2(_10388_),
    .B1(\line_cache[86][4] ),
    .B2(_10389_),
    .C1(_11343_),
    .X(_11344_));
 sky130_fd_sc_hd__a22o_1 _15623_ (.A1(_10396_),
    .A2(\line_cache[88][4] ),
    .B1(_10397_),
    .B2(\line_cache[89][4] ),
    .X(_11345_));
 sky130_fd_sc_hd__a221o_1 _15624_ (.A1(\line_cache[91][4] ),
    .A2(_10394_),
    .B1(\line_cache[90][4] ),
    .B2(_10395_),
    .C1(_11345_),
    .X(_11346_));
 sky130_fd_sc_hd__or4_1 _15625_ (.A(_11340_),
    .B(_11342_),
    .C(_11344_),
    .D(_11346_),
    .X(_11347_));
 sky130_fd_sc_hd__a22o_1 _15626_ (.A1(_10371_),
    .A2(\line_cache[100][4] ),
    .B1(_10372_),
    .B2(\line_cache[101][4] ),
    .X(_11348_));
 sky130_fd_sc_hd__a22o_1 _15627_ (.A1(_10369_),
    .A2(\line_cache[103][4] ),
    .B1(_10370_),
    .B2(\line_cache[102][4] ),
    .X(_11349_));
 sky130_fd_sc_hd__a22o_1 _15628_ (.A1(_10351_),
    .A2(\line_cache[96][4] ),
    .B1(_10352_),
    .B2(\line_cache[97][4] ),
    .X(_11350_));
 sky130_fd_sc_hd__a221o_2 _15629_ (.A1(\line_cache[99][4] ),
    .A2(_10349_),
    .B1(\line_cache[98][4] ),
    .B2(_10348_),
    .C1(_11350_),
    .X(_11351_));
 sky130_fd_sc_hd__and3_1 _15630_ (.A(_10035_),
    .B(\line_cache[107][4] ),
    .C(_10651_),
    .X(_11352_));
 sky130_fd_sc_hd__and3_1 _15631_ (.A(_10176_),
    .B(\line_cache[105][4] ),
    .C(_10651_),
    .X(_11353_));
 sky130_fd_sc_hd__and3_1 _15632_ (.A(_10054_),
    .B(\line_cache[106][4] ),
    .C(_10356_),
    .X(_11354_));
 sky130_fd_sc_hd__and3_1 _15633_ (.A(_10360_),
    .B(\line_cache[104][4] ),
    .C(_10356_),
    .X(_11355_));
 sky130_fd_sc_hd__or4_1 _15634_ (.A(_11352_),
    .B(_11353_),
    .C(_11354_),
    .D(_11355_),
    .X(_11356_));
 sky130_fd_sc_hd__a22o_1 _15635_ (.A1(_10365_),
    .A2(\line_cache[108][4] ),
    .B1(_10366_),
    .B2(\line_cache[109][4] ),
    .X(_11357_));
 sky130_fd_sc_hd__a221o_1 _15636_ (.A1(\line_cache[111][4] ),
    .A2(_10363_),
    .B1(\line_cache[110][4] ),
    .B2(_10364_),
    .C1(_11357_),
    .X(_11358_));
 sky130_fd_sc_hd__or2_1 _15637_ (.A(_11356_),
    .B(_11358_),
    .X(_11359_));
 sky130_fd_sc_hd__or4_1 _15638_ (.A(_11348_),
    .B(_11349_),
    .C(_11351_),
    .D(_11359_),
    .X(_11360_));
 sky130_fd_sc_hd__nor2_1 _15639_ (.A(_11347_),
    .B(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__and3_1 _15640_ (.A(_10176_),
    .B(\line_cache[121][4] ),
    .C(_10302_),
    .X(_11362_));
 sky130_fd_sc_hd__a21o_1 _15641_ (.A1(\line_cache[120][4] ),
    .A2(_10317_),
    .B1(_11362_),
    .X(_11363_));
 sky130_fd_sc_hd__a221o_1 _15642_ (.A1(\line_cache[123][4] ),
    .A2(_10315_),
    .B1(\line_cache[122][4] ),
    .B2(_10316_),
    .C1(_11363_),
    .X(_11364_));
 sky130_fd_sc_hd__a22o_1 _15643_ (.A1(_10298_),
    .A2(\line_cache[112][4] ),
    .B1(_10299_),
    .B2(\line_cache[113][4] ),
    .X(_11365_));
 sky130_fd_sc_hd__a221o_1 _15644_ (.A1(\line_cache[115][4] ),
    .A2(_10296_),
    .B1(\line_cache[114][4] ),
    .B2(_10297_),
    .C1(_11365_),
    .X(_11366_));
 sky130_fd_sc_hd__a22o_1 _15645_ (.A1(_10311_),
    .A2(\line_cache[116][4] ),
    .B1(_10312_),
    .B2(\line_cache[117][4] ),
    .X(_11367_));
 sky130_fd_sc_hd__a221o_1 _15646_ (.A1(\line_cache[119][4] ),
    .A2(_10309_),
    .B1(\line_cache[118][4] ),
    .B2(_10310_),
    .C1(_11367_),
    .X(_11368_));
 sky130_fd_sc_hd__a22o_1 _15647_ (.A1(_10305_),
    .A2(\line_cache[124][4] ),
    .B1(_10306_),
    .B2(\line_cache[125][4] ),
    .X(_11369_));
 sky130_fd_sc_hd__a221o_1 _15648_ (.A1(\line_cache[126][4] ),
    .A2(_10304_),
    .B1(\line_cache[127][4] ),
    .B2(_10622_),
    .C1(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__or4_1 _15649_ (.A(_11364_),
    .B(_11366_),
    .C(_11368_),
    .D(_11370_),
    .X(_11371_));
 sky130_fd_sc_hd__and3_1 _15650_ (.A(_09758_),
    .B(_10098_),
    .C(\line_cache[133][4] ),
    .X(_11372_));
 sky130_fd_sc_hd__a21o_1 _15651_ (.A1(\line_cache[132][4] ),
    .A2(_10324_),
    .B1(_11372_),
    .X(_11373_));
 sky130_fd_sc_hd__a221o_1 _15652_ (.A1(\line_cache[135][4] ),
    .A2(_10322_),
    .B1(\line_cache[134][4] ),
    .B2(_10323_),
    .C1(_11373_),
    .X(_11374_));
 sky130_fd_sc_hd__a22o_1 _15653_ (.A1(_10330_),
    .A2(\line_cache[129][4] ),
    .B1(\line_cache[128][4] ),
    .B2(_10629_),
    .X(_11375_));
 sky130_fd_sc_hd__a221o_1 _15654_ (.A1(\line_cache[131][4] ),
    .A2(_10328_),
    .B1(\line_cache[130][4] ),
    .B2(_10329_),
    .C1(_11375_),
    .X(_11376_));
 sky130_fd_sc_hd__a22o_1 _15655_ (.A1(_10342_),
    .A2(\line_cache[139][4] ),
    .B1(\line_cache[138][4] ),
    .B2(_10343_),
    .X(_11377_));
 sky130_fd_sc_hd__a221o_1 _15656_ (.A1(\line_cache[137][4] ),
    .A2(_10340_),
    .B1(\line_cache[136][4] ),
    .B2(_10341_),
    .C1(_11377_),
    .X(_11378_));
 sky130_fd_sc_hd__a22o_1 _15657_ (.A1(_10336_),
    .A2(\line_cache[140][4] ),
    .B1(\line_cache[141][4] ),
    .B2(_10337_),
    .X(_11379_));
 sky130_fd_sc_hd__a221o_1 _15658_ (.A1(\line_cache[143][4] ),
    .A2(_10334_),
    .B1(\line_cache[142][4] ),
    .B2(_10335_),
    .C1(_11379_),
    .X(_11380_));
 sky130_fd_sc_hd__or4_2 _15659_ (.A(_11374_),
    .B(_11376_),
    .C(_11378_),
    .D(_11380_),
    .X(_11381_));
 sky130_fd_sc_hd__nor2_1 _15660_ (.A(_11371_),
    .B(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__a22o_1 _15661_ (.A1(_10244_),
    .A2(\line_cache[173][4] ),
    .B1(\line_cache[172][4] ),
    .B2(_10245_),
    .X(_11383_));
 sky130_fd_sc_hd__a221o_1 _15662_ (.A1(\line_cache[175][4] ),
    .A2(_10242_),
    .B1(\line_cache[174][4] ),
    .B2(_10243_),
    .C1(_11383_),
    .X(_11384_));
 sky130_fd_sc_hd__a22o_1 _15663_ (.A1(_10250_),
    .A2(\line_cache[165][4] ),
    .B1(\line_cache[164][4] ),
    .B2(_10251_),
    .X(_11385_));
 sky130_fd_sc_hd__a221oi_1 _15664_ (.A1(\line_cache[167][4] ),
    .A2(_10248_),
    .B1(\line_cache[166][4] ),
    .B2(_10249_),
    .C1(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__a22o_1 _15665_ (.A1(_10256_),
    .A2(\line_cache[160][4] ),
    .B1(\line_cache[161][4] ),
    .B2(_10257_),
    .X(_11387_));
 sky130_fd_sc_hd__a221oi_4 _15666_ (.A1(\line_cache[163][4] ),
    .A2(_10254_),
    .B1(\line_cache[162][4] ),
    .B2(_10255_),
    .C1(_11387_),
    .Y(_11388_));
 sky130_fd_sc_hd__a22o_1 _15667_ (.A1(_10261_),
    .A2(\line_cache[168][4] ),
    .B1(\line_cache[169][4] ),
    .B2(_10260_),
    .X(_11389_));
 sky130_fd_sc_hd__a221oi_2 _15668_ (.A1(\line_cache[171][4] ),
    .A2(_10262_),
    .B1(\line_cache[170][4] ),
    .B2(_10263_),
    .C1(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__and4b_1 _15669_ (.A_N(_11384_),
    .B(_11386_),
    .C(_11388_),
    .D(_11390_),
    .X(_11391_));
 sky130_fd_sc_hd__a22o_1 _15670_ (.A1(_10277_),
    .A2(\line_cache[184][4] ),
    .B1(\line_cache[185][4] ),
    .B2(_10278_),
    .X(_11392_));
 sky130_fd_sc_hd__a221o_1 _15671_ (.A1(\line_cache[187][4] ),
    .A2(_10275_),
    .B1(\line_cache[186][4] ),
    .B2(_10276_),
    .C1(_11392_),
    .X(_11393_));
 sky130_fd_sc_hd__a22o_1 _15672_ (.A1(_10284_),
    .A2(\line_cache[176][4] ),
    .B1(_10285_),
    .B2(\line_cache[177][4] ),
    .X(_11394_));
 sky130_fd_sc_hd__a221oi_2 _15673_ (.A1(\line_cache[179][4] ),
    .A2(_10282_),
    .B1(\line_cache[178][4] ),
    .B2(_10283_),
    .C1(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__and3_1 _15674_ (.A(_10288_),
    .B(_10102_),
    .C(\line_cache[182][4] ),
    .X(_11396_));
 sky130_fd_sc_hd__and3_1 _15675_ (.A(_10288_),
    .B(_10098_),
    .C(\line_cache[181][4] ),
    .X(_11397_));
 sky130_fd_sc_hd__a31o_1 _15676_ (.A1(\line_cache[180][4] ),
    .A2(_10288_),
    .A3(_10106_),
    .B1(_11397_),
    .X(_11398_));
 sky130_fd_sc_hd__a311oi_2 _15677_ (.A1(\line_cache[183][4] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_11396_),
    .C1(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__a22o_1 _15678_ (.A1(_10272_),
    .A2(\line_cache[189][4] ),
    .B1(\line_cache[188][4] ),
    .B2(_10271_),
    .X(_11400_));
 sky130_fd_sc_hd__a221oi_1 _15679_ (.A1(\line_cache[191][4] ),
    .A2(_10269_),
    .B1(\line_cache[190][4] ),
    .B2(_10270_),
    .C1(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__and4b_1 _15680_ (.A_N(_11393_),
    .B(_11395_),
    .C(_11399_),
    .D(_11401_),
    .X(_11402_));
 sky130_fd_sc_hd__a22o_1 _15681_ (.A1(_10219_),
    .A2(\line_cache[157][4] ),
    .B1(\line_cache[156][4] ),
    .B2(_10220_),
    .X(_11403_));
 sky130_fd_sc_hd__a221o_1 _15682_ (.A1(\line_cache[159][4] ),
    .A2(_10217_),
    .B1(\line_cache[158][4] ),
    .B2(_10218_),
    .C1(_11403_),
    .X(_11404_));
 sky130_fd_sc_hd__a22o_1 _15683_ (.A1(_10238_),
    .A2(\line_cache[154][4] ),
    .B1(\line_cache[155][4] ),
    .B2(_10237_),
    .X(_11405_));
 sky130_fd_sc_hd__a221o_1 _15684_ (.A1(\line_cache[153][4] ),
    .A2(_10235_),
    .B1(\line_cache[152][4] ),
    .B2(_10236_),
    .C1(_11405_),
    .X(_11406_));
 sky130_fd_sc_hd__a22o_1 _15685_ (.A1(_10224_),
    .A2(\line_cache[148][4] ),
    .B1(\line_cache[149][4] ),
    .B2(_10223_),
    .X(_11407_));
 sky130_fd_sc_hd__a22o_1 _15686_ (.A1(_10225_),
    .A2(\line_cache[151][4] ),
    .B1(\line_cache[150][4] ),
    .B2(_10226_),
    .X(_11408_));
 sky130_fd_sc_hd__a22o_1 _15687_ (.A1(_10230_),
    .A2(\line_cache[144][4] ),
    .B1(\line_cache[145][4] ),
    .B2(_10229_),
    .X(_11409_));
 sky130_fd_sc_hd__a22o_1 _15688_ (.A1(_10231_),
    .A2(\line_cache[147][4] ),
    .B1(\line_cache[146][4] ),
    .B2(_10232_),
    .X(_11410_));
 sky130_fd_sc_hd__or4_1 _15689_ (.A(_11407_),
    .B(_11408_),
    .C(_11409_),
    .D(_11410_),
    .X(_11411_));
 sky130_fd_sc_hd__nor3_1 _15690_ (.A(_11404_),
    .B(_11406_),
    .C(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__and3_2 _15691_ (.A(_11391_),
    .B(_11402_),
    .C(_11412_),
    .X(_11413_));
 sky130_fd_sc_hd__and3_1 _15692_ (.A(_11361_),
    .B(_11382_),
    .C(_11413_),
    .X(_11414_));
 sky130_fd_sc_hd__nand3_1 _15693_ (.A(_11275_),
    .B(_11338_),
    .C(_11414_),
    .Y(_11415_));
 sky130_fd_sc_hd__o21ba_2 _15694_ (.A1(_11168_),
    .A2(_11415_),
    .B1_N(_08979_),
    .X(_11416_));
 sky130_fd_sc_hd__buf_6 _15695_ (.A(_11416_),
    .X(net130));
 sky130_fd_sc_hd__and2_1 _15696_ (.A(_09912_),
    .B(\line_cache[0][5] ),
    .X(_11417_));
 sky130_fd_sc_hd__and3_1 _15697_ (.A(_10102_),
    .B(\line_cache[70][5] ),
    .C(_10161_),
    .X(_11418_));
 sky130_fd_sc_hd__a22o_1 _15698_ (.A1(_10163_),
    .A2(\line_cache[68][5] ),
    .B1(_10164_),
    .B2(\line_cache[69][5] ),
    .X(_11419_));
 sky130_fd_sc_hd__a211o_1 _15699_ (.A1(\line_cache[71][5] ),
    .A2(_10159_),
    .B1(_11418_),
    .C1(_11419_),
    .X(_11420_));
 sky130_fd_sc_hd__and3_1 _15700_ (.A(_10031_),
    .B(\line_cache[77][5] ),
    .C(_10167_),
    .X(_11421_));
 sky130_fd_sc_hd__and3_1 _15701_ (.A(_10038_),
    .B(\line_cache[78][5] ),
    .C(_10167_),
    .X(_11422_));
 sky130_fd_sc_hd__and3_1 _15702_ (.A(_10041_),
    .B(\line_cache[76][5] ),
    .C(_10161_),
    .X(_11423_));
 sky130_fd_sc_hd__a2111o_1 _15703_ (.A1(_10168_),
    .A2(\line_cache[79][5] ),
    .B1(_11421_),
    .C1(_11422_),
    .D1(_11423_),
    .X(_11424_));
 sky130_fd_sc_hd__and3_1 _15704_ (.A(_10176_),
    .B(\line_cache[73][5] ),
    .C(_10160_),
    .X(_11425_));
 sky130_fd_sc_hd__a21o_1 _15705_ (.A1(\line_cache[72][5] ),
    .A2(_10175_),
    .B1(_11425_),
    .X(_11426_));
 sky130_fd_sc_hd__a221o_1 _15706_ (.A1(\line_cache[75][5] ),
    .A2(_10173_),
    .B1(\line_cache[74][5] ),
    .B2(_10174_),
    .C1(_11426_),
    .X(_11427_));
 sky130_fd_sc_hd__a22o_1 _15707_ (.A1(_10182_),
    .A2(\line_cache[64][5] ),
    .B1(_10183_),
    .B2(\line_cache[65][5] ),
    .X(_11428_));
 sky130_fd_sc_hd__a221o_1 _15708_ (.A1(\line_cache[67][5] ),
    .A2(_10180_),
    .B1(\line_cache[66][5] ),
    .B2(_10181_),
    .C1(_11428_),
    .X(_11429_));
 sky130_fd_sc_hd__or4_2 _15709_ (.A(_11420_),
    .B(_11424_),
    .C(_11427_),
    .D(_11429_),
    .X(_11430_));
 sky130_fd_sc_hd__a22o_1 _15710_ (.A1(_10189_),
    .A2(\line_cache[252][5] ),
    .B1(_10190_),
    .B2(\line_cache[251][5] ),
    .X(_11431_));
 sky130_fd_sc_hd__a221o_1 _15711_ (.A1(\line_cache[254][5] ),
    .A2(_10187_),
    .B1(\line_cache[253][5] ),
    .B2(_10188_),
    .C1(_11431_),
    .X(_11432_));
 sky130_fd_sc_hd__a22o_1 _15712_ (.A1(_10195_),
    .A2(\line_cache[248][5] ),
    .B1(_10196_),
    .B2(\line_cache[247][5] ),
    .X(_11433_));
 sky130_fd_sc_hd__a221o_1 _15713_ (.A1(\line_cache[250][5] ),
    .A2(_10193_),
    .B1(\line_cache[249][5] ),
    .B2(_10194_),
    .C1(_11433_),
    .X(_11434_));
 sky130_fd_sc_hd__and2b_1 _15714_ (.A_N(_10200_),
    .B(\line_cache[240][5] ),
    .X(_11435_));
 sky130_fd_sc_hd__and2b_1 _15715_ (.A_N(_09570_),
    .B(\line_cache[241][5] ),
    .X(_11436_));
 sky130_fd_sc_hd__and2b_1 _15716_ (.A_N(_10203_),
    .B(\line_cache[242][5] ),
    .X(_11437_));
 sky130_fd_sc_hd__a2111o_1 _15717_ (.A1(\line_cache[239][5] ),
    .A2(_10199_),
    .B1(_11435_),
    .C1(_11436_),
    .D1(_11437_),
    .X(_11438_));
 sky130_fd_sc_hd__and2b_1 _15718_ (.A_N(_10206_),
    .B(\line_cache[243][5] ),
    .X(_11439_));
 sky130_fd_sc_hd__and2b_1 _15719_ (.A_N(_10208_),
    .B(\line_cache[244][5] ),
    .X(_11440_));
 sky130_fd_sc_hd__and2b_1 _15720_ (.A_N(_09597_),
    .B(\line_cache[245][5] ),
    .X(_11441_));
 sky130_fd_sc_hd__and2b_1 _15721_ (.A_N(_10211_),
    .B(\line_cache[246][5] ),
    .X(_11442_));
 sky130_fd_sc_hd__or4_1 _15722_ (.A(_11439_),
    .B(_11440_),
    .C(_11441_),
    .D(_11442_),
    .X(_11443_));
 sky130_fd_sc_hd__or4_1 _15723_ (.A(_11432_),
    .B(_11434_),
    .C(_11438_),
    .D(_11443_),
    .X(_11444_));
 sky130_fd_sc_hd__and3_1 _15724_ (.A(_09595_),
    .B(\line_cache[229][5] ),
    .C(_10099_),
    .X(_11445_));
 sky130_fd_sc_hd__and3_1 _15725_ (.A(_10044_),
    .B(\line_cache[230][5] ),
    .C(_10099_),
    .X(_11446_));
 sky130_fd_sc_hd__and3_1 _15726_ (.A(_10104_),
    .B(\line_cache[227][5] ),
    .C(_10434_),
    .X(_11447_));
 sky130_fd_sc_hd__and3_1 _15727_ (.A(_10106_),
    .B(\line_cache[228][5] ),
    .C(_10437_),
    .X(_11448_));
 sky130_fd_sc_hd__or4_1 _15728_ (.A(_11445_),
    .B(_11446_),
    .C(_11447_),
    .D(_11448_),
    .X(_11449_));
 sky130_fd_sc_hd__and3_1 _15729_ (.A(_09544_),
    .B(\line_cache[223][5] ),
    .C(_10109_),
    .X(_11450_));
 sky130_fd_sc_hd__and3_1 _15730_ (.A(_10070_),
    .B(\line_cache[224][5] ),
    .C(_10434_),
    .X(_11451_));
 sky130_fd_sc_hd__and3_1 _15731_ (.A(_10067_),
    .B(\line_cache[225][5] ),
    .C(_10437_),
    .X(_11452_));
 sky130_fd_sc_hd__and3_1 _15732_ (.A(_10074_),
    .B(\line_cache[226][5] ),
    .C(_10437_),
    .X(_11453_));
 sky130_fd_sc_hd__or4_1 _15733_ (.A(_11450_),
    .B(_11451_),
    .C(_11452_),
    .D(_11453_),
    .X(_11454_));
 sky130_fd_sc_hd__a22o_1 _15734_ (.A1(_10118_),
    .A2(\line_cache[236][5] ),
    .B1(_10120_),
    .B2(\line_cache[235][5] ),
    .X(_11455_));
 sky130_fd_sc_hd__a221o_1 _15735_ (.A1(\line_cache[238][5] ),
    .A2(_10116_),
    .B1(\line_cache[237][5] ),
    .B2(_10117_),
    .C1(_11455_),
    .X(_11456_));
 sky130_fd_sc_hd__a22o_1 _15736_ (.A1(_10125_),
    .A2(\line_cache[232][5] ),
    .B1(_10126_),
    .B2(\line_cache[231][5] ),
    .X(_11457_));
 sky130_fd_sc_hd__a221o_1 _15737_ (.A1(\line_cache[234][5] ),
    .A2(_10123_),
    .B1(\line_cache[233][5] ),
    .B2(_10124_),
    .C1(_11457_),
    .X(_11458_));
 sky130_fd_sc_hd__or4_1 _15738_ (.A(_11449_),
    .B(_11454_),
    .C(_11456_),
    .D(_11458_),
    .X(_11459_));
 sky130_fd_sc_hd__a22o_1 _15739_ (.A1(_10132_),
    .A2(\line_cache[220][5] ),
    .B1(_10133_),
    .B2(\line_cache[219][5] ),
    .X(_11460_));
 sky130_fd_sc_hd__a221o_1 _15740_ (.A1(\line_cache[222][5] ),
    .A2(_10130_),
    .B1(\line_cache[221][5] ),
    .B2(_10131_),
    .C1(_11460_),
    .X(_11461_));
 sky130_fd_sc_hd__a22o_1 _15741_ (.A1(_10138_),
    .A2(\line_cache[208][5] ),
    .B1(_10139_),
    .B2(\line_cache[207][5] ),
    .X(_11462_));
 sky130_fd_sc_hd__a221o_1 _15742_ (.A1(\line_cache[210][5] ),
    .A2(_10136_),
    .B1(\line_cache[209][5] ),
    .B2(_10137_),
    .C1(_11462_),
    .X(_11463_));
 sky130_fd_sc_hd__a22o_1 _15743_ (.A1(_10144_),
    .A2(\line_cache[216][5] ),
    .B1(_10145_),
    .B2(\line_cache[215][5] ),
    .X(_11464_));
 sky130_fd_sc_hd__a221o_1 _15744_ (.A1(\line_cache[218][5] ),
    .A2(_10142_),
    .B1(\line_cache[217][5] ),
    .B2(_10143_),
    .C1(_11464_),
    .X(_11465_));
 sky130_fd_sc_hd__and2b_1 _15745_ (.A_N(_10148_),
    .B(\line_cache[211][5] ),
    .X(_11466_));
 sky130_fd_sc_hd__nor2b_1 _15746_ (.A(_10150_),
    .B_N(\line_cache[212][5] ),
    .Y(_11467_));
 sky130_fd_sc_hd__and2b_1 _15747_ (.A_N(_10152_),
    .B(\line_cache[213][5] ),
    .X(_11468_));
 sky130_fd_sc_hd__and2b_1 _15748_ (.A_N(_10154_),
    .B(\line_cache[214][5] ),
    .X(_11469_));
 sky130_fd_sc_hd__or4_1 _15749_ (.A(_11466_),
    .B(_11467_),
    .C(_11468_),
    .D(_11469_),
    .X(_11470_));
 sky130_fd_sc_hd__or4_2 _15750_ (.A(_11461_),
    .B(_11463_),
    .C(_11465_),
    .D(_11470_),
    .X(_11471_));
 sky130_fd_sc_hd__or2_1 _15751_ (.A(_11459_),
    .B(_11471_),
    .X(_11472_));
 sky130_fd_sc_hd__or3_1 _15752_ (.A(_11430_),
    .B(_11444_),
    .C(_11472_),
    .X(_11473_));
 sky130_fd_sc_hd__and3_1 _15753_ (.A(_10035_),
    .B(\line_cache[203][5] ),
    .C(_09539_),
    .X(_11474_));
 sky130_fd_sc_hd__and3_1 _15754_ (.A(_10038_),
    .B(\line_cache[206][5] ),
    .C(_10075_),
    .X(_11475_));
 sky130_fd_sc_hd__and3_1 _15755_ (.A(_10041_),
    .B(\line_cache[204][5] ),
    .C(_10075_),
    .X(_11476_));
 sky130_fd_sc_hd__a2111o_1 _15756_ (.A1(\line_cache[205][5] ),
    .A2(_10033_),
    .B1(_11474_),
    .C1(_11475_),
    .D1(_11476_),
    .X(_11477_));
 sky130_fd_sc_hd__a22o_1 _15757_ (.A1(_10049_),
    .A2(\line_cache[195][5] ),
    .B1(\line_cache[196][5] ),
    .B2(_10051_),
    .X(_11478_));
 sky130_fd_sc_hd__a221o_1 _15758_ (.A1(\line_cache[198][5] ),
    .A2(_10046_),
    .B1(\line_cache[197][5] ),
    .B2(_10047_),
    .C1(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__a22o_1 _15759_ (.A1(_10060_),
    .A2(\line_cache[200][5] ),
    .B1(_10063_),
    .B2(\line_cache[199][5] ),
    .X(_11480_));
 sky130_fd_sc_hd__a221o_1 _15760_ (.A1(\line_cache[202][5] ),
    .A2(_10056_),
    .B1(\line_cache[201][5] ),
    .B2(_10059_),
    .C1(_11480_),
    .X(_11481_));
 sky130_fd_sc_hd__and3_1 _15761_ (.A(_10067_),
    .B(\line_cache[193][5] ),
    .C(_10075_),
    .X(_11482_));
 sky130_fd_sc_hd__and3_1 _15762_ (.A(_10071_),
    .B(\line_cache[192][5] ),
    .C(_09540_),
    .X(_11483_));
 sky130_fd_sc_hd__and3_1 _15763_ (.A(_10074_),
    .B(\line_cache[194][5] ),
    .C(_09540_),
    .X(_11484_));
 sky130_fd_sc_hd__a2111o_1 _15764_ (.A1(_10066_),
    .A2(\line_cache[286][5] ),
    .B1(_11482_),
    .C1(_11483_),
    .D1(_11484_),
    .X(_11485_));
 sky130_fd_sc_hd__or4_1 _15765_ (.A(_11477_),
    .B(_11479_),
    .C(_11481_),
    .D(_11485_),
    .X(_11486_));
 sky130_fd_sc_hd__a22o_1 _15766_ (.A1(_09623_),
    .A2(\line_cache[275][5] ),
    .B1(_09620_),
    .B2(\line_cache[274][5] ),
    .X(_11487_));
 sky130_fd_sc_hd__a22o_1 _15767_ (.A1(_10080_),
    .A2(\line_cache[276][5] ),
    .B1(\line_cache[277][5] ),
    .B2(_10081_),
    .X(_11488_));
 sky130_fd_sc_hd__a22o_1 _15768_ (.A1(_10086_),
    .A2(\line_cache[270][5] ),
    .B1(\line_cache[269][5] ),
    .B2(_10088_),
    .X(_11489_));
 sky130_fd_sc_hd__a221o_1 _15769_ (.A1(\line_cache[273][5] ),
    .A2(_10083_),
    .B1(\line_cache[272][5] ),
    .B2(_10084_),
    .C1(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__a22o_1 _15770_ (.A1(_09658_),
    .A2(\line_cache[283][5] ),
    .B1(\line_cache[282][5] ),
    .B2(_09661_),
    .X(_11491_));
 sky130_fd_sc_hd__a22o_1 _15771_ (.A1(_09645_),
    .A2(\line_cache[285][5] ),
    .B1(\line_cache[284][5] ),
    .B2(_09648_),
    .X(_11492_));
 sky130_fd_sc_hd__a22o_1 _15772_ (.A1(_09639_),
    .A2(\line_cache[279][5] ),
    .B1(\line_cache[278][5] ),
    .B2(_09636_),
    .X(_11493_));
 sky130_fd_sc_hd__a221o_1 _15773_ (.A1(\line_cache[281][5] ),
    .A2(_09663_),
    .B1(\line_cache[280][5] ),
    .B2(_09655_),
    .C1(_11493_),
    .X(_11494_));
 sky130_fd_sc_hd__or3_1 _15774_ (.A(_11491_),
    .B(_11492_),
    .C(_11494_),
    .X(_11495_));
 sky130_fd_sc_hd__or4_1 _15775_ (.A(_11487_),
    .B(_11488_),
    .C(_11490_),
    .D(_11495_),
    .X(_11496_));
 sky130_fd_sc_hd__nor2_1 _15776_ (.A(_11486_),
    .B(_11496_),
    .Y(_11497_));
 sky130_fd_sc_hd__and2b_1 _15777_ (.A_N(_09987_),
    .B(\line_cache[256][5] ),
    .X(_11498_));
 sky130_fd_sc_hd__and2b_1 _15778_ (.A_N(_09747_),
    .B(\line_cache[302][5] ),
    .X(_11499_));
 sky130_fd_sc_hd__a22o_1 _15779_ (.A1(_09743_),
    .A2(\line_cache[301][5] ),
    .B1(\line_cache[300][5] ),
    .B2(_09742_),
    .X(_11500_));
 sky130_fd_sc_hd__or3_1 _15780_ (.A(_11498_),
    .B(_11499_),
    .C(_11500_),
    .X(_11501_));
 sky130_fd_sc_hd__and3_1 _15781_ (.A(_09917_),
    .B(_09691_),
    .C(\line_cache[258][5] ),
    .X(_11502_));
 sky130_fd_sc_hd__and3_1 _15782_ (.A(_09848_),
    .B(_09691_),
    .C(\line_cache[260][5] ),
    .X(_11503_));
 sky130_fd_sc_hd__and3_1 _15783_ (.A(_09919_),
    .B(_09611_),
    .C(\line_cache[257][5] ),
    .X(_11504_));
 sky130_fd_sc_hd__and3_1 _15784_ (.A(_09840_),
    .B(_09611_),
    .C(\line_cache[259][5] ),
    .X(_11505_));
 sky130_fd_sc_hd__or4_1 _15785_ (.A(_11502_),
    .B(_11503_),
    .C(_11504_),
    .D(_11505_),
    .X(_11506_));
 sky130_fd_sc_hd__and3_1 _15786_ (.A(_09858_),
    .B(_09547_),
    .C(\line_cache[267][5] ),
    .X(_11507_));
 sky130_fd_sc_hd__a22o_1 _15787_ (.A1(_09998_),
    .A2(\line_cache[265][5] ),
    .B1(\line_cache[266][5] ),
    .B2(_09999_),
    .X(_11508_));
 sky130_fd_sc_hd__a311o_1 _15788_ (.A1(_09548_),
    .A2(\line_cache[268][5] ),
    .A3(_09862_),
    .B1(_11507_),
    .C1(_11508_),
    .X(_11509_));
 sky130_fd_sc_hd__nand2_1 _15789_ (.A(_10007_),
    .B(\line_cache[262][5] ),
    .Y(_11510_));
 sky130_fd_sc_hd__nand2_1 _15790_ (.A(_10010_),
    .B(\line_cache[261][5] ),
    .Y(_11511_));
 sky130_fd_sc_hd__nand2_1 _15791_ (.A(_11510_),
    .B(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__a221oi_1 _15792_ (.A1(_10003_),
    .A2(\line_cache[264][5] ),
    .B1(_10005_),
    .B2(\line_cache[263][5] ),
    .C1(_11512_),
    .Y(_11513_));
 sky130_fd_sc_hd__or4b_1 _15793_ (.A(_11501_),
    .B(_11506_),
    .C(_11509_),
    .D_N(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__a22o_1 _15794_ (.A1(_09682_),
    .A2(\line_cache[308][5] ),
    .B1(\line_cache[309][5] ),
    .B2(_09685_),
    .X(_11515_));
 sky130_fd_sc_hd__a221o_1 _15795_ (.A1(\line_cache[311][5] ),
    .A2(_09689_),
    .B1(\line_cache[310][5] ),
    .B2(_09693_),
    .C1(_11515_),
    .X(_11516_));
 sky130_fd_sc_hd__a22o_1 _15796_ (.A1(_09728_),
    .A2(\line_cache[295][5] ),
    .B1(\line_cache[294][5] ),
    .B2(_09726_),
    .X(_11517_));
 sky130_fd_sc_hd__a221o_1 _15797_ (.A1(\line_cache[293][5] ),
    .A2(_09730_),
    .B1(\line_cache[292][5] ),
    .B2(_10018_),
    .C1(_11517_),
    .X(_11518_));
 sky130_fd_sc_hd__a22o_1 _15798_ (.A1(_09716_),
    .A2(\line_cache[296][5] ),
    .B1(\line_cache[297][5] ),
    .B2(_09721_),
    .X(_11519_));
 sky130_fd_sc_hd__a221o_1 _15799_ (.A1(\line_cache[299][5] ),
    .A2(_09718_),
    .B1(\line_cache[298][5] ),
    .B2(_09720_),
    .C1(_11519_),
    .X(_11520_));
 sky130_fd_sc_hd__a22o_1 _15800_ (.A1(_10025_),
    .A2(\line_cache[288][5] ),
    .B1(\line_cache[289][5] ),
    .B2(_10026_),
    .X(_11521_));
 sky130_fd_sc_hd__a221o_1 _15801_ (.A1(\line_cache[291][5] ),
    .A2(_10023_),
    .B1(\line_cache[290][5] ),
    .B2(_10024_),
    .C1(_11521_),
    .X(_11522_));
 sky130_fd_sc_hd__or4_2 _15802_ (.A(_11516_),
    .B(_11518_),
    .C(_11520_),
    .D(_11522_),
    .X(_11523_));
 sky130_fd_sc_hd__nor2_1 _15803_ (.A(_11514_),
    .B(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__nand2_1 _15804_ (.A(_11497_),
    .B(_11524_),
    .Y(_11525_));
 sky130_fd_sc_hd__nor2_1 _15805_ (.A(_11473_),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__a22o_1 _15806_ (.A1(_09842_),
    .A2(\line_cache[6][5] ),
    .B1(\line_cache[5][5] ),
    .B2(_09844_),
    .X(_11527_));
 sky130_fd_sc_hd__a221o_1 _15807_ (.A1(\line_cache[4][5] ),
    .A2(_09850_),
    .B1(\line_cache[3][5] ),
    .B2(_09914_),
    .C1(_11527_),
    .X(_11528_));
 sky130_fd_sc_hd__and3_1 _15808_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][5] ),
    .X(_11529_));
 sky130_fd_sc_hd__and3_1 _15809_ (.A(_09919_),
    .B(_09533_),
    .C(\line_cache[1][5] ),
    .X(_11530_));
 sky130_fd_sc_hd__a211o_1 _15810_ (.A1(\line_cache[15][5] ),
    .A2(_09867_),
    .B1(_11529_),
    .C1(_11530_),
    .X(_11531_));
 sky130_fd_sc_hd__and3_1 _15811_ (.A(_09922_),
    .B(_09531_),
    .C(\line_cache[63][5] ),
    .X(_11532_));
 sky130_fd_sc_hd__a31o_1 _15812_ (.A1(_09547_),
    .A2(\line_cache[319][5] ),
    .A3(_09922_),
    .B1(_11532_),
    .X(_11533_));
 sky130_fd_sc_hd__a221o_1 _15813_ (.A1(\line_cache[47][5] ),
    .A2(_09806_),
    .B1(\line_cache[31][5] ),
    .B2(_09907_),
    .C1(_11533_),
    .X(_11534_));
 sky130_fd_sc_hd__nand2_1 _15814_ (.A(_09746_),
    .B(\line_cache[303][5] ),
    .Y(_11535_));
 sky130_fd_sc_hd__nand2_1 _15815_ (.A(_09930_),
    .B(\line_cache[271][5] ),
    .Y(_11536_));
 sky130_fd_sc_hd__nand2_1 _15816_ (.A(_11535_),
    .B(_11536_),
    .Y(_11537_));
 sky130_fd_sc_hd__a221oi_2 _15817_ (.A1(\line_cache[255][5] ),
    .A2(_09926_),
    .B1(\line_cache[287][5] ),
    .B2(_09927_),
    .C1(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__or4b_1 _15818_ (.A(_11528_),
    .B(_11531_),
    .C(_11534_),
    .D_N(_11538_),
    .X(_11539_));
 sky130_fd_sc_hd__a22o_1 _15819_ (.A1(_09803_),
    .A2(\line_cache[45][5] ),
    .B1(\line_cache[46][5] ),
    .B2(_09804_),
    .X(_11540_));
 sky130_fd_sc_hd__a22o_1 _15820_ (.A1(_09824_),
    .A2(\line_cache[48][5] ),
    .B1(\line_cache[49][5] ),
    .B2(_09826_),
    .X(_11541_));
 sky130_fd_sc_hd__nand2_1 _15821_ (.A(_09787_),
    .B(\line_cache[41][5] ),
    .Y(_11542_));
 sky130_fd_sc_hd__nand2_1 _15822_ (.A(_09789_),
    .B(\line_cache[42][5] ),
    .Y(_11543_));
 sky130_fd_sc_hd__nand2_1 _15823_ (.A(_11542_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__a221oi_2 _15824_ (.A1(_09785_),
    .A2(\line_cache[43][5] ),
    .B1(\line_cache[44][5] ),
    .B2(_09801_),
    .C1(_11544_),
    .Y(_11545_));
 sky130_fd_sc_hd__or3b_1 _15825_ (.A(_11540_),
    .B(_11541_),
    .C_N(_11545_),
    .X(_11546_));
 sky130_fd_sc_hd__a22o_1 _15826_ (.A1(_09699_),
    .A2(\line_cache[317][5] ),
    .B1(\line_cache[316][5] ),
    .B2(_09697_),
    .X(_11547_));
 sky130_fd_sc_hd__a22o_1 _15827_ (.A1(_09832_),
    .A2(\line_cache[58][5] ),
    .B1(\line_cache[59][5] ),
    .B2(_09833_),
    .X(_11548_));
 sky130_fd_sc_hd__a22o_1 _15828_ (.A1(_09819_),
    .A2(\line_cache[61][5] ),
    .B1(\line_cache[60][5] ),
    .B2(_09817_),
    .X(_11549_));
 sky130_fd_sc_hd__a22o_1 _15829_ (.A1(_09822_),
    .A2(\line_cache[62][5] ),
    .B1(\line_cache[318][5] ),
    .B2(_09702_),
    .X(_11550_));
 sky130_fd_sc_hd__or4_1 _15830_ (.A(_11547_),
    .B(_11548_),
    .C(_11549_),
    .D(_11550_),
    .X(_11551_));
 sky130_fd_sc_hd__a22o_1 _15831_ (.A1(_09675_),
    .A2(\line_cache[304][5] ),
    .B1(\line_cache[305][5] ),
    .B2(_09676_),
    .X(_11552_));
 sky130_fd_sc_hd__a22o_1 _15832_ (.A1(_09705_),
    .A2(\line_cache[312][5] ),
    .B1(\line_cache[313][5] ),
    .B2(_09707_),
    .X(_11553_));
 sky130_fd_sc_hd__a22o_1 _15833_ (.A1(_09708_),
    .A2(\line_cache[314][5] ),
    .B1(\line_cache[315][5] ),
    .B2(_09709_),
    .X(_11554_));
 sky130_fd_sc_hd__a22o_1 _15834_ (.A1(_09677_),
    .A2(\line_cache[306][5] ),
    .B1(\line_cache[307][5] ),
    .B2(_09678_),
    .X(_11555_));
 sky130_fd_sc_hd__or4_1 _15835_ (.A(_11552_),
    .B(_11553_),
    .C(_11554_),
    .D(_11555_),
    .X(_11556_));
 sky130_fd_sc_hd__a22o_1 _15836_ (.A1(_09830_),
    .A2(\line_cache[56][5] ),
    .B1(\line_cache[57][5] ),
    .B2(_09834_),
    .X(_11557_));
 sky130_fd_sc_hd__a22o_1 _15837_ (.A1(_09809_),
    .A2(\line_cache[52][5] ),
    .B1(\line_cache[53][5] ),
    .B2(_09811_),
    .X(_11558_));
 sky130_fd_sc_hd__a22o_1 _15838_ (.A1(_09827_),
    .A2(\line_cache[50][5] ),
    .B1(\line_cache[51][5] ),
    .B2(_09828_),
    .X(_11559_));
 sky130_fd_sc_hd__a22o_1 _15839_ (.A1(_09813_),
    .A2(\line_cache[54][5] ),
    .B1(\line_cache[55][5] ),
    .B2(_09815_),
    .X(_11560_));
 sky130_fd_sc_hd__or4_1 _15840_ (.A(_11557_),
    .B(_11558_),
    .C(_11559_),
    .D(_11560_),
    .X(_11561_));
 sky130_fd_sc_hd__or4_2 _15841_ (.A(_11546_),
    .B(_11551_),
    .C(_11556_),
    .D(_11561_),
    .X(_11562_));
 sky130_fd_sc_hd__nand2_1 _15842_ (.A(_09864_),
    .B(\line_cache[12][5] ),
    .Y(_11563_));
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(_09860_),
    .B(\line_cache[11][5] ),
    .Y(_11564_));
 sky130_fd_sc_hd__nand2_1 _15844_ (.A(_11563_),
    .B(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__a221oi_2 _15845_ (.A1(_09870_),
    .A2(\line_cache[14][5] ),
    .B1(\line_cache[13][5] ),
    .B2(_09873_),
    .C1(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__nand2_1 _15846_ (.A(_09853_),
    .B(\line_cache[10][5] ),
    .Y(_11567_));
 sky130_fd_sc_hd__nand2_1 _15847_ (.A(_09857_),
    .B(\line_cache[9][5] ),
    .Y(_11568_));
 sky130_fd_sc_hd__nand2_1 _15848_ (.A(_11567_),
    .B(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__a221oi_1 _15849_ (.A1(_09855_),
    .A2(\line_cache[8][5] ),
    .B1(_09847_),
    .B2(\line_cache[7][5] ),
    .C1(_11569_),
    .Y(_11570_));
 sky130_fd_sc_hd__nand2_1 _15850_ (.A(_11566_),
    .B(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__and3_1 _15851_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][5] ),
    .X(_11572_));
 sky130_fd_sc_hd__a22o_1 _15852_ (.A1(_09884_),
    .A2(\line_cache[23][5] ),
    .B1(\line_cache[22][5] ),
    .B2(_09886_),
    .X(_11573_));
 sky130_fd_sc_hd__a22o_1 _15853_ (.A1(_09877_),
    .A2(\line_cache[19][5] ),
    .B1(\line_cache[18][5] ),
    .B2(_09878_),
    .X(_11574_));
 sky130_fd_sc_hd__a221o_1 _15854_ (.A1(\line_cache[17][5] ),
    .A2(_09969_),
    .B1(\line_cache[16][5] ),
    .B2(_09970_),
    .C1(_11574_),
    .X(_11575_));
 sky130_fd_sc_hd__a2111o_1 _15855_ (.A1(\line_cache[20][5] ),
    .A2(_09888_),
    .B1(_11572_),
    .C1(_11573_),
    .D1(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__a22o_1 _15856_ (.A1(_09796_),
    .A2(\line_cache[33][5] ),
    .B1(\line_cache[34][5] ),
    .B2(_09798_),
    .X(_11577_));
 sky130_fd_sc_hd__a221o_1 _15857_ (.A1(\line_cache[36][5] ),
    .A2(_09777_),
    .B1(\line_cache[35][5] ),
    .B2(_09794_),
    .C1(_11577_),
    .X(_11578_));
 sky130_fd_sc_hd__a22o_1 _15858_ (.A1(_09890_),
    .A2(\line_cache[27][5] ),
    .B1(\line_cache[26][5] ),
    .B2(_09896_),
    .X(_11579_));
 sky130_fd_sc_hd__a221oi_2 _15859_ (.A1(\line_cache[25][5] ),
    .A2(_09892_),
    .B1(\line_cache[24][5] ),
    .B2(_09895_),
    .C1(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__a22o_1 _15860_ (.A1(_09903_),
    .A2(\line_cache[29][5] ),
    .B1(\line_cache[28][5] ),
    .B2(_09900_),
    .X(_11581_));
 sky130_fd_sc_hd__a221oi_1 _15861_ (.A1(\line_cache[32][5] ),
    .A2(_09792_),
    .B1(\line_cache[30][5] ),
    .B2(_09905_),
    .C1(_11581_),
    .Y(_11582_));
 sky130_fd_sc_hd__nand2_1 _15862_ (.A(_09773_),
    .B(\line_cache[38][5] ),
    .Y(_11583_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_09775_),
    .B(\line_cache[37][5] ),
    .Y(_11584_));
 sky130_fd_sc_hd__nand2_1 _15864_ (.A(_11583_),
    .B(_11584_),
    .Y(_11585_));
 sky130_fd_sc_hd__a221oi_2 _15865_ (.A1(_09783_),
    .A2(\line_cache[40][5] ),
    .B1(\line_cache[39][5] ),
    .B2(_09780_),
    .C1(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__and4b_1 _15866_ (.A_N(_11578_),
    .B(_11580_),
    .C(_11582_),
    .D(_11586_),
    .X(_11587_));
 sky130_fd_sc_hd__or3b_1 _15867_ (.A(_11571_),
    .B(_11576_),
    .C_N(_11587_),
    .X(_11588_));
 sky130_fd_sc_hd__nor3_2 _15868_ (.A(_11539_),
    .B(_11562_),
    .C(_11588_),
    .Y(_11589_));
 sky130_fd_sc_hd__a22o_1 _15869_ (.A1(_10219_),
    .A2(\line_cache[157][5] ),
    .B1(\line_cache[156][5] ),
    .B2(_10220_),
    .X(_11590_));
 sky130_fd_sc_hd__a221o_1 _15870_ (.A1(\line_cache[159][5] ),
    .A2(_10217_),
    .B1(\line_cache[158][5] ),
    .B2(_10218_),
    .C1(_11590_),
    .X(_11591_));
 sky130_fd_sc_hd__a22o_1 _15871_ (.A1(_10238_),
    .A2(\line_cache[154][5] ),
    .B1(\line_cache[155][5] ),
    .B2(_10237_),
    .X(_11592_));
 sky130_fd_sc_hd__a221o_1 _15872_ (.A1(\line_cache[153][5] ),
    .A2(_10235_),
    .B1(\line_cache[152][5] ),
    .B2(_10236_),
    .C1(_11592_),
    .X(_11593_));
 sky130_fd_sc_hd__and4_1 _15873_ (.A(_09753_),
    .B(_09532_),
    .C(\line_cache[149][5] ),
    .D(_09683_),
    .X(_11594_));
 sky130_fd_sc_hd__a22o_1 _15874_ (.A1(_10225_),
    .A2(\line_cache[151][5] ),
    .B1(\line_cache[150][5] ),
    .B2(_10226_),
    .X(_11595_));
 sky130_fd_sc_hd__a22o_1 _15875_ (.A1(_10230_),
    .A2(\line_cache[144][5] ),
    .B1(\line_cache[145][5] ),
    .B2(_10229_),
    .X(_11596_));
 sky130_fd_sc_hd__a221o_1 _15876_ (.A1(\line_cache[147][5] ),
    .A2(_10231_),
    .B1(\line_cache[146][5] ),
    .B2(_10232_),
    .C1(_11596_),
    .X(_11597_));
 sky130_fd_sc_hd__a2111o_1 _15877_ (.A1(\line_cache[148][5] ),
    .A2(_10224_),
    .B1(_11594_),
    .C1(_11595_),
    .D1(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__nor3_1 _15878_ (.A(_11591_),
    .B(_11593_),
    .C(_11598_),
    .Y(_11599_));
 sky130_fd_sc_hd__a22o_1 _15879_ (.A1(_10277_),
    .A2(\line_cache[184][5] ),
    .B1(\line_cache[185][5] ),
    .B2(_10278_),
    .X(_11600_));
 sky130_fd_sc_hd__a221o_1 _15880_ (.A1(\line_cache[187][5] ),
    .A2(_10275_),
    .B1(\line_cache[186][5] ),
    .B2(_10276_),
    .C1(_11600_),
    .X(_11601_));
 sky130_fd_sc_hd__a22o_1 _15881_ (.A1(_10284_),
    .A2(\line_cache[176][5] ),
    .B1(_10285_),
    .B2(\line_cache[177][5] ),
    .X(_11602_));
 sky130_fd_sc_hd__a221oi_2 _15882_ (.A1(\line_cache[179][5] ),
    .A2(_10282_),
    .B1(\line_cache[178][5] ),
    .B2(_10283_),
    .C1(_11602_),
    .Y(_11603_));
 sky130_fd_sc_hd__and3_1 _15883_ (.A(_10288_),
    .B(_10102_),
    .C(\line_cache[182][5] ),
    .X(_11604_));
 sky130_fd_sc_hd__and3_1 _15884_ (.A(_10288_),
    .B(_10098_),
    .C(\line_cache[181][5] ),
    .X(_11605_));
 sky130_fd_sc_hd__a31o_1 _15885_ (.A1(\line_cache[180][5] ),
    .A2(_10289_),
    .A3(_10106_),
    .B1(_11605_),
    .X(_11606_));
 sky130_fd_sc_hd__a311oi_2 _15886_ (.A1(\line_cache[183][5] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_11604_),
    .C1(_11606_),
    .Y(_11607_));
 sky130_fd_sc_hd__a22o_1 _15887_ (.A1(_10272_),
    .A2(\line_cache[189][5] ),
    .B1(\line_cache[188][5] ),
    .B2(_10271_),
    .X(_11608_));
 sky130_fd_sc_hd__a221oi_1 _15888_ (.A1(\line_cache[191][5] ),
    .A2(_10269_),
    .B1(\line_cache[190][5] ),
    .B2(_10270_),
    .C1(_11608_),
    .Y(_11609_));
 sky130_fd_sc_hd__and4b_1 _15889_ (.A_N(_11601_),
    .B(_11603_),
    .C(_11607_),
    .D(_11609_),
    .X(_11610_));
 sky130_fd_sc_hd__a22o_1 _15890_ (.A1(_10244_),
    .A2(\line_cache[173][5] ),
    .B1(\line_cache[172][5] ),
    .B2(_10245_),
    .X(_11611_));
 sky130_fd_sc_hd__a221o_1 _15891_ (.A1(\line_cache[175][5] ),
    .A2(_10242_),
    .B1(\line_cache[174][5] ),
    .B2(_10243_),
    .C1(_11611_),
    .X(_11612_));
 sky130_fd_sc_hd__a22o_1 _15892_ (.A1(_10263_),
    .A2(\line_cache[170][5] ),
    .B1(\line_cache[171][5] ),
    .B2(_10262_),
    .X(_11613_));
 sky130_fd_sc_hd__a221o_1 _15893_ (.A1(\line_cache[169][5] ),
    .A2(_10260_),
    .B1(\line_cache[168][5] ),
    .B2(_10261_),
    .C1(_11613_),
    .X(_11614_));
 sky130_fd_sc_hd__a22o_1 _15894_ (.A1(_10256_),
    .A2(\line_cache[160][5] ),
    .B1(\line_cache[161][5] ),
    .B2(_10257_),
    .X(_11615_));
 sky130_fd_sc_hd__a22o_1 _15895_ (.A1(_10250_),
    .A2(\line_cache[165][5] ),
    .B1(\line_cache[164][5] ),
    .B2(_10251_),
    .X(_11616_));
 sky130_fd_sc_hd__a22o_1 _15896_ (.A1(_10248_),
    .A2(\line_cache[167][5] ),
    .B1(\line_cache[166][5] ),
    .B2(_10249_),
    .X(_11617_));
 sky130_fd_sc_hd__a22o_1 _15897_ (.A1(_10255_),
    .A2(\line_cache[162][5] ),
    .B1(\line_cache[163][5] ),
    .B2(_10254_),
    .X(_11618_));
 sky130_fd_sc_hd__or4_1 _15898_ (.A(_11615_),
    .B(_11616_),
    .C(_11617_),
    .D(_11618_),
    .X(_11619_));
 sky130_fd_sc_hd__nor3_1 _15899_ (.A(_11612_),
    .B(_11614_),
    .C(_11619_),
    .Y(_11620_));
 sky130_fd_sc_hd__and3_2 _15900_ (.A(_11599_),
    .B(_11610_),
    .C(_11620_),
    .X(_11621_));
 sky130_fd_sc_hd__a22o_1 _15901_ (.A1(_10378_),
    .A2(\line_cache[80][5] ),
    .B1(_10379_),
    .B2(\line_cache[81][5] ),
    .X(_11622_));
 sky130_fd_sc_hd__a221o_1 _15902_ (.A1(\line_cache[83][5] ),
    .A2(_10376_),
    .B1(\line_cache[82][5] ),
    .B2(_10377_),
    .C1(_11622_),
    .X(_11623_));
 sky130_fd_sc_hd__a22o_1 _15903_ (.A1(_10384_),
    .A2(\line_cache[92][5] ),
    .B1(_10385_),
    .B2(\line_cache[93][5] ),
    .X(_11624_));
 sky130_fd_sc_hd__a221o_1 _15904_ (.A1(\line_cache[95][5] ),
    .A2(net136),
    .B1(\line_cache[94][5] ),
    .B2(_10383_),
    .C1(_11624_),
    .X(_11625_));
 sky130_fd_sc_hd__a22o_1 _15905_ (.A1(_10390_),
    .A2(\line_cache[84][5] ),
    .B1(_10391_),
    .B2(\line_cache[85][5] ),
    .X(_11626_));
 sky130_fd_sc_hd__a221o_1 _15906_ (.A1(\line_cache[87][5] ),
    .A2(_10388_),
    .B1(\line_cache[86][5] ),
    .B2(_10389_),
    .C1(_11626_),
    .X(_11627_));
 sky130_fd_sc_hd__a22o_1 _15907_ (.A1(_10396_),
    .A2(\line_cache[88][5] ),
    .B1(_10397_),
    .B2(\line_cache[89][5] ),
    .X(_11628_));
 sky130_fd_sc_hd__a221o_1 _15908_ (.A1(\line_cache[91][5] ),
    .A2(_10394_),
    .B1(\line_cache[90][5] ),
    .B2(_10395_),
    .C1(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__or4_1 _15909_ (.A(_11623_),
    .B(_11625_),
    .C(_11627_),
    .D(_11629_),
    .X(_11630_));
 sky130_fd_sc_hd__a22o_1 _15910_ (.A1(_10371_),
    .A2(\line_cache[100][5] ),
    .B1(_10372_),
    .B2(\line_cache[101][5] ),
    .X(_11631_));
 sky130_fd_sc_hd__a22o_1 _15911_ (.A1(_10369_),
    .A2(\line_cache[103][5] ),
    .B1(_10370_),
    .B2(\line_cache[102][5] ),
    .X(_11632_));
 sky130_fd_sc_hd__a22o_1 _15912_ (.A1(_10351_),
    .A2(\line_cache[96][5] ),
    .B1(_10352_),
    .B2(\line_cache[97][5] ),
    .X(_11633_));
 sky130_fd_sc_hd__a221o_2 _15913_ (.A1(\line_cache[99][5] ),
    .A2(_10349_),
    .B1(\line_cache[98][5] ),
    .B2(_10348_),
    .C1(_11633_),
    .X(_11634_));
 sky130_fd_sc_hd__and3_1 _15914_ (.A(_10035_),
    .B(\line_cache[107][5] ),
    .C(_10651_),
    .X(_11635_));
 sky130_fd_sc_hd__and3_1 _15915_ (.A(_10176_),
    .B(\line_cache[105][5] ),
    .C(_10651_),
    .X(_11636_));
 sky130_fd_sc_hd__and3_1 _15916_ (.A(_10054_),
    .B(\line_cache[106][5] ),
    .C(_10356_),
    .X(_11637_));
 sky130_fd_sc_hd__and3_1 _15917_ (.A(_10360_),
    .B(\line_cache[104][5] ),
    .C(_10356_),
    .X(_11638_));
 sky130_fd_sc_hd__or4_1 _15918_ (.A(_11635_),
    .B(_11636_),
    .C(_11637_),
    .D(_11638_),
    .X(_11639_));
 sky130_fd_sc_hd__a22o_1 _15919_ (.A1(_10365_),
    .A2(\line_cache[108][5] ),
    .B1(_10366_),
    .B2(\line_cache[109][5] ),
    .X(_11640_));
 sky130_fd_sc_hd__a221o_1 _15920_ (.A1(\line_cache[111][5] ),
    .A2(_10363_),
    .B1(\line_cache[110][5] ),
    .B2(_10364_),
    .C1(_11640_),
    .X(_11641_));
 sky130_fd_sc_hd__or2_1 _15921_ (.A(_11639_),
    .B(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__or4_1 _15922_ (.A(_11631_),
    .B(_11632_),
    .C(_11634_),
    .D(_11642_),
    .X(_11643_));
 sky130_fd_sc_hd__nor2_1 _15923_ (.A(_11630_),
    .B(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__and3_1 _15924_ (.A(_10176_),
    .B(\line_cache[121][5] ),
    .C(_10302_),
    .X(_11645_));
 sky130_fd_sc_hd__a21o_1 _15925_ (.A1(\line_cache[120][5] ),
    .A2(_10317_),
    .B1(_11645_),
    .X(_11646_));
 sky130_fd_sc_hd__a221o_1 _15926_ (.A1(\line_cache[123][5] ),
    .A2(_10315_),
    .B1(\line_cache[122][5] ),
    .B2(_10316_),
    .C1(_11646_),
    .X(_11647_));
 sky130_fd_sc_hd__a22o_1 _15927_ (.A1(_10298_),
    .A2(\line_cache[112][5] ),
    .B1(_10299_),
    .B2(\line_cache[113][5] ),
    .X(_11648_));
 sky130_fd_sc_hd__a221o_1 _15928_ (.A1(\line_cache[115][5] ),
    .A2(_10296_),
    .B1(\line_cache[114][5] ),
    .B2(_10297_),
    .C1(_11648_),
    .X(_11649_));
 sky130_fd_sc_hd__a22o_1 _15929_ (.A1(_10311_),
    .A2(\line_cache[116][5] ),
    .B1(_10312_),
    .B2(\line_cache[117][5] ),
    .X(_11650_));
 sky130_fd_sc_hd__a221o_1 _15930_ (.A1(\line_cache[119][5] ),
    .A2(_10309_),
    .B1(\line_cache[118][5] ),
    .B2(_10310_),
    .C1(_11650_),
    .X(_11651_));
 sky130_fd_sc_hd__a22o_1 _15931_ (.A1(_10305_),
    .A2(\line_cache[124][5] ),
    .B1(_10306_),
    .B2(\line_cache[125][5] ),
    .X(_11652_));
 sky130_fd_sc_hd__a221o_1 _15932_ (.A1(\line_cache[126][5] ),
    .A2(_10304_),
    .B1(\line_cache[127][5] ),
    .B2(_10622_),
    .C1(_11652_),
    .X(_11653_));
 sky130_fd_sc_hd__or4_1 _15933_ (.A(_11647_),
    .B(_11649_),
    .C(_11651_),
    .D(_11653_),
    .X(_11654_));
 sky130_fd_sc_hd__a22o_1 _15934_ (.A1(_10322_),
    .A2(\line_cache[135][5] ),
    .B1(\line_cache[134][5] ),
    .B2(_10323_),
    .X(_11655_));
 sky130_fd_sc_hd__a221o_1 _15935_ (.A1(\line_cache[133][5] ),
    .A2(_10626_),
    .B1(\line_cache[132][5] ),
    .B2(_10324_),
    .C1(_11655_),
    .X(_11656_));
 sky130_fd_sc_hd__a22o_1 _15936_ (.A1(_10330_),
    .A2(\line_cache[129][5] ),
    .B1(\line_cache[128][5] ),
    .B2(_10629_),
    .X(_11657_));
 sky130_fd_sc_hd__a221o_1 _15937_ (.A1(\line_cache[131][5] ),
    .A2(_10328_),
    .B1(\line_cache[130][5] ),
    .B2(_10329_),
    .C1(_11657_),
    .X(_11658_));
 sky130_fd_sc_hd__a22o_1 _15938_ (.A1(_10336_),
    .A2(\line_cache[140][5] ),
    .B1(\line_cache[141][5] ),
    .B2(_10337_),
    .X(_11659_));
 sky130_fd_sc_hd__a221o_1 _15939_ (.A1(\line_cache[143][5] ),
    .A2(_10334_),
    .B1(\line_cache[142][5] ),
    .B2(_10335_),
    .C1(_11659_),
    .X(_11660_));
 sky130_fd_sc_hd__a22o_1 _15940_ (.A1(_10342_),
    .A2(\line_cache[139][5] ),
    .B1(\line_cache[138][5] ),
    .B2(_10343_),
    .X(_11661_));
 sky130_fd_sc_hd__a221o_1 _15941_ (.A1(\line_cache[137][5] ),
    .A2(_10340_),
    .B1(\line_cache[136][5] ),
    .B2(_10341_),
    .C1(_11661_),
    .X(_11662_));
 sky130_fd_sc_hd__or4_2 _15942_ (.A(_11656_),
    .B(_11658_),
    .C(_11660_),
    .D(_11662_),
    .X(_11663_));
 sky130_fd_sc_hd__nor2_1 _15943_ (.A(_11654_),
    .B(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__and3_1 _15944_ (.A(_11621_),
    .B(_11644_),
    .C(_11664_),
    .X(_11665_));
 sky130_fd_sc_hd__nand3_1 _15945_ (.A(_11526_),
    .B(_11589_),
    .C(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__o21ba_2 _15946_ (.A1(_11417_),
    .A2(_11666_),
    .B1_N(_08979_),
    .X(_11667_));
 sky130_fd_sc_hd__buf_6 _15947_ (.A(_11667_),
    .X(net131));
 sky130_fd_sc_hd__and2_1 _15948_ (.A(_09912_),
    .B(\line_cache[0][6] ),
    .X(_11668_));
 sky130_fd_sc_hd__and3_1 _15949_ (.A(_10031_),
    .B(\line_cache[77][6] ),
    .C(_10167_),
    .X(_11669_));
 sky130_fd_sc_hd__and3_1 _15950_ (.A(_10038_),
    .B(\line_cache[78][6] ),
    .C(_10167_),
    .X(_11670_));
 sky130_fd_sc_hd__and3_1 _15951_ (.A(_10041_),
    .B(\line_cache[76][6] ),
    .C(_10161_),
    .X(_11671_));
 sky130_fd_sc_hd__a2111o_1 _15952_ (.A1(_10168_),
    .A2(\line_cache[79][6] ),
    .B1(_11669_),
    .C1(_11670_),
    .D1(_11671_),
    .X(_11672_));
 sky130_fd_sc_hd__a22o_1 _15953_ (.A1(_10182_),
    .A2(\line_cache[64][6] ),
    .B1(_10183_),
    .B2(\line_cache[65][6] ),
    .X(_11673_));
 sky130_fd_sc_hd__a221o_1 _15954_ (.A1(\line_cache[67][6] ),
    .A2(_10180_),
    .B1(\line_cache[66][6] ),
    .B2(_10181_),
    .C1(_11673_),
    .X(_11674_));
 sky130_fd_sc_hd__a22o_1 _15955_ (.A1(_10163_),
    .A2(\line_cache[68][6] ),
    .B1(_10164_),
    .B2(\line_cache[69][6] ),
    .X(_11675_));
 sky130_fd_sc_hd__a221o_1 _15956_ (.A1(\line_cache[71][6] ),
    .A2(_10159_),
    .B1(\line_cache[70][6] ),
    .B2(_10750_),
    .C1(_11675_),
    .X(_11676_));
 sky130_fd_sc_hd__a22o_1 _15957_ (.A1(_10175_),
    .A2(\line_cache[72][6] ),
    .B1(_10753_),
    .B2(\line_cache[73][6] ),
    .X(_11677_));
 sky130_fd_sc_hd__a221o_1 _15958_ (.A1(\line_cache[75][6] ),
    .A2(_10173_),
    .B1(\line_cache[74][6] ),
    .B2(_10174_),
    .C1(_11677_),
    .X(_11678_));
 sky130_fd_sc_hd__or4_4 _15959_ (.A(_11672_),
    .B(_11674_),
    .C(_11676_),
    .D(_11678_),
    .X(_11679_));
 sky130_fd_sc_hd__a22o_1 _15960_ (.A1(_10189_),
    .A2(\line_cache[252][6] ),
    .B1(_10190_),
    .B2(\line_cache[251][6] ),
    .X(_11680_));
 sky130_fd_sc_hd__a221o_1 _15961_ (.A1(\line_cache[254][6] ),
    .A2(_10187_),
    .B1(\line_cache[253][6] ),
    .B2(_10188_),
    .C1(_11680_),
    .X(_11681_));
 sky130_fd_sc_hd__a22o_1 _15962_ (.A1(_10195_),
    .A2(\line_cache[248][6] ),
    .B1(_10196_),
    .B2(\line_cache[247][6] ),
    .X(_11682_));
 sky130_fd_sc_hd__a221o_1 _15963_ (.A1(\line_cache[250][6] ),
    .A2(_10193_),
    .B1(\line_cache[249][6] ),
    .B2(_10194_),
    .C1(_11682_),
    .X(_11683_));
 sky130_fd_sc_hd__and2b_1 _15964_ (.A_N(_10200_),
    .B(\line_cache[240][6] ),
    .X(_11684_));
 sky130_fd_sc_hd__and2b_1 _15965_ (.A_N(_09570_),
    .B(\line_cache[241][6] ),
    .X(_11685_));
 sky130_fd_sc_hd__and2b_1 _15966_ (.A_N(_10203_),
    .B(\line_cache[242][6] ),
    .X(_11686_));
 sky130_fd_sc_hd__a2111o_1 _15967_ (.A1(\line_cache[239][6] ),
    .A2(_10199_),
    .B1(_11684_),
    .C1(_11685_),
    .D1(_11686_),
    .X(_11687_));
 sky130_fd_sc_hd__and2b_1 _15968_ (.A_N(_10206_),
    .B(\line_cache[243][6] ),
    .X(_11688_));
 sky130_fd_sc_hd__and2b_1 _15969_ (.A_N(_10208_),
    .B(\line_cache[244][6] ),
    .X(_11689_));
 sky130_fd_sc_hd__and2b_1 _15970_ (.A_N(_09597_),
    .B(\line_cache[245][6] ),
    .X(_11690_));
 sky130_fd_sc_hd__and2b_1 _15971_ (.A_N(_10211_),
    .B(\line_cache[246][6] ),
    .X(_11691_));
 sky130_fd_sc_hd__or4_1 _15972_ (.A(_11688_),
    .B(_11689_),
    .C(_11690_),
    .D(_11691_),
    .X(_11692_));
 sky130_fd_sc_hd__or4_1 _15973_ (.A(_11681_),
    .B(_11683_),
    .C(_11687_),
    .D(_11692_),
    .X(_11693_));
 sky130_fd_sc_hd__and3_1 _15974_ (.A(_09595_),
    .B(\line_cache[229][6] ),
    .C(_10099_),
    .X(_11694_));
 sky130_fd_sc_hd__and3_1 _15975_ (.A(_10044_),
    .B(\line_cache[230][6] ),
    .C(_10099_),
    .X(_11695_));
 sky130_fd_sc_hd__and3_1 _15976_ (.A(_10104_),
    .B(\line_cache[227][6] ),
    .C(_10434_),
    .X(_11696_));
 sky130_fd_sc_hd__and3_1 _15977_ (.A(_10106_),
    .B(\line_cache[228][6] ),
    .C(_10437_),
    .X(_11697_));
 sky130_fd_sc_hd__or4_1 _15978_ (.A(_11694_),
    .B(_11695_),
    .C(_11696_),
    .D(_11697_),
    .X(_11698_));
 sky130_fd_sc_hd__and3_1 _15979_ (.A(_09544_),
    .B(\line_cache[223][6] ),
    .C(_10109_),
    .X(_11699_));
 sky130_fd_sc_hd__and3_1 _15980_ (.A(_10070_),
    .B(\line_cache[224][6] ),
    .C(_10434_),
    .X(_11700_));
 sky130_fd_sc_hd__and3_1 _15981_ (.A(_10067_),
    .B(\line_cache[225][6] ),
    .C(_10437_),
    .X(_11701_));
 sky130_fd_sc_hd__and3_1 _15982_ (.A(_10074_),
    .B(\line_cache[226][6] ),
    .C(_10437_),
    .X(_11702_));
 sky130_fd_sc_hd__or4_1 _15983_ (.A(_11699_),
    .B(_11700_),
    .C(_11701_),
    .D(_11702_),
    .X(_11703_));
 sky130_fd_sc_hd__a22o_1 _15984_ (.A1(_10118_),
    .A2(\line_cache[236][6] ),
    .B1(_10120_),
    .B2(\line_cache[235][6] ),
    .X(_11704_));
 sky130_fd_sc_hd__a221o_1 _15985_ (.A1(\line_cache[238][6] ),
    .A2(_10116_),
    .B1(\line_cache[237][6] ),
    .B2(_10117_),
    .C1(_11704_),
    .X(_11705_));
 sky130_fd_sc_hd__a22o_1 _15986_ (.A1(_10125_),
    .A2(\line_cache[232][6] ),
    .B1(_10126_),
    .B2(\line_cache[231][6] ),
    .X(_11706_));
 sky130_fd_sc_hd__a221o_1 _15987_ (.A1(\line_cache[234][6] ),
    .A2(_10123_),
    .B1(\line_cache[233][6] ),
    .B2(_10124_),
    .C1(_11706_),
    .X(_11707_));
 sky130_fd_sc_hd__or4_1 _15988_ (.A(_11698_),
    .B(_11703_),
    .C(_11705_),
    .D(_11707_),
    .X(_11708_));
 sky130_fd_sc_hd__a22o_1 _15989_ (.A1(_10132_),
    .A2(\line_cache[220][6] ),
    .B1(_10133_),
    .B2(\line_cache[219][6] ),
    .X(_11709_));
 sky130_fd_sc_hd__a221o_1 _15990_ (.A1(\line_cache[222][6] ),
    .A2(_10130_),
    .B1(\line_cache[221][6] ),
    .B2(_10131_),
    .C1(_11709_),
    .X(_11710_));
 sky130_fd_sc_hd__a22o_1 _15991_ (.A1(_10138_),
    .A2(\line_cache[208][6] ),
    .B1(_10139_),
    .B2(\line_cache[207][6] ),
    .X(_11711_));
 sky130_fd_sc_hd__a221o_1 _15992_ (.A1(\line_cache[210][6] ),
    .A2(_10136_),
    .B1(\line_cache[209][6] ),
    .B2(_10137_),
    .C1(_11711_),
    .X(_11712_));
 sky130_fd_sc_hd__a22o_1 _15993_ (.A1(_10144_),
    .A2(\line_cache[216][6] ),
    .B1(_10145_),
    .B2(\line_cache[215][6] ),
    .X(_11713_));
 sky130_fd_sc_hd__a221o_1 _15994_ (.A1(\line_cache[218][6] ),
    .A2(_10142_),
    .B1(\line_cache[217][6] ),
    .B2(_10143_),
    .C1(_11713_),
    .X(_11714_));
 sky130_fd_sc_hd__and2b_1 _15995_ (.A_N(_10148_),
    .B(\line_cache[211][6] ),
    .X(_11715_));
 sky130_fd_sc_hd__nor2b_1 _15996_ (.A(_10150_),
    .B_N(\line_cache[212][6] ),
    .Y(_11716_));
 sky130_fd_sc_hd__and2b_1 _15997_ (.A_N(_10152_),
    .B(\line_cache[213][6] ),
    .X(_11717_));
 sky130_fd_sc_hd__and2b_1 _15998_ (.A_N(_10154_),
    .B(\line_cache[214][6] ),
    .X(_11718_));
 sky130_fd_sc_hd__or4_1 _15999_ (.A(_11715_),
    .B(_11716_),
    .C(_11717_),
    .D(_11718_),
    .X(_11719_));
 sky130_fd_sc_hd__or4_2 _16000_ (.A(_11710_),
    .B(_11712_),
    .C(_11714_),
    .D(_11719_),
    .X(_11720_));
 sky130_fd_sc_hd__or2_1 _16001_ (.A(_11708_),
    .B(_11720_),
    .X(_11721_));
 sky130_fd_sc_hd__or3_1 _16002_ (.A(_11679_),
    .B(_11693_),
    .C(_11721_),
    .X(_11722_));
 sky130_fd_sc_hd__and3_1 _16003_ (.A(_10035_),
    .B(\line_cache[203][6] ),
    .C(_09539_),
    .X(_11723_));
 sky130_fd_sc_hd__and3_1 _16004_ (.A(_10038_),
    .B(\line_cache[206][6] ),
    .C(_10075_),
    .X(_11724_));
 sky130_fd_sc_hd__and3_1 _16005_ (.A(_10041_),
    .B(\line_cache[204][6] ),
    .C(_10075_),
    .X(_11725_));
 sky130_fd_sc_hd__a2111o_1 _16006_ (.A1(\line_cache[205][6] ),
    .A2(_10033_),
    .B1(_11723_),
    .C1(_11724_),
    .D1(_11725_),
    .X(_11726_));
 sky130_fd_sc_hd__a22o_1 _16007_ (.A1(_10049_),
    .A2(\line_cache[195][6] ),
    .B1(\line_cache[196][6] ),
    .B2(_10051_),
    .X(_11727_));
 sky130_fd_sc_hd__a221o_1 _16008_ (.A1(\line_cache[198][6] ),
    .A2(_10046_),
    .B1(\line_cache[197][6] ),
    .B2(_10047_),
    .C1(_11727_),
    .X(_11728_));
 sky130_fd_sc_hd__a22o_1 _16009_ (.A1(_10060_),
    .A2(\line_cache[200][6] ),
    .B1(_10063_),
    .B2(\line_cache[199][6] ),
    .X(_11729_));
 sky130_fd_sc_hd__a221o_1 _16010_ (.A1(\line_cache[202][6] ),
    .A2(_10056_),
    .B1(\line_cache[201][6] ),
    .B2(_10059_),
    .C1(_11729_),
    .X(_11730_));
 sky130_fd_sc_hd__and3_1 _16011_ (.A(_10067_),
    .B(\line_cache[193][6] ),
    .C(_10075_),
    .X(_11731_));
 sky130_fd_sc_hd__and3_1 _16012_ (.A(_10071_),
    .B(\line_cache[192][6] ),
    .C(_09540_),
    .X(_11732_));
 sky130_fd_sc_hd__and3_1 _16013_ (.A(_10074_),
    .B(\line_cache[194][6] ),
    .C(_09540_),
    .X(_11733_));
 sky130_fd_sc_hd__a2111o_1 _16014_ (.A1(_10066_),
    .A2(\line_cache[286][6] ),
    .B1(_11731_),
    .C1(_11732_),
    .D1(_11733_),
    .X(_11734_));
 sky130_fd_sc_hd__or4_2 _16015_ (.A(_11726_),
    .B(_11728_),
    .C(_11730_),
    .D(_11734_),
    .X(_11735_));
 sky130_fd_sc_hd__a22o_1 _16016_ (.A1(_09623_),
    .A2(\line_cache[275][6] ),
    .B1(_09620_),
    .B2(\line_cache[274][6] ),
    .X(_11736_));
 sky130_fd_sc_hd__a22o_1 _16017_ (.A1(_10080_),
    .A2(\line_cache[276][6] ),
    .B1(\line_cache[277][6] ),
    .B2(_10081_),
    .X(_11737_));
 sky130_fd_sc_hd__a22o_1 _16018_ (.A1(_10086_),
    .A2(\line_cache[270][6] ),
    .B1(\line_cache[269][6] ),
    .B2(_10088_),
    .X(_11738_));
 sky130_fd_sc_hd__a221o_1 _16019_ (.A1(\line_cache[273][6] ),
    .A2(_10083_),
    .B1(\line_cache[272][6] ),
    .B2(_10084_),
    .C1(_11738_),
    .X(_11739_));
 sky130_fd_sc_hd__a22o_1 _16020_ (.A1(_09658_),
    .A2(\line_cache[283][6] ),
    .B1(\line_cache[282][6] ),
    .B2(_09661_),
    .X(_11740_));
 sky130_fd_sc_hd__a22o_1 _16021_ (.A1(_09645_),
    .A2(\line_cache[285][6] ),
    .B1(\line_cache[284][6] ),
    .B2(_09648_),
    .X(_11741_));
 sky130_fd_sc_hd__a22o_1 _16022_ (.A1(_09639_),
    .A2(\line_cache[279][6] ),
    .B1(\line_cache[278][6] ),
    .B2(_09636_),
    .X(_11742_));
 sky130_fd_sc_hd__a221o_1 _16023_ (.A1(\line_cache[281][6] ),
    .A2(_09663_),
    .B1(\line_cache[280][6] ),
    .B2(_09655_),
    .C1(_11742_),
    .X(_11743_));
 sky130_fd_sc_hd__or3_1 _16024_ (.A(_11740_),
    .B(_11741_),
    .C(_11743_),
    .X(_11744_));
 sky130_fd_sc_hd__or4_1 _16025_ (.A(_11736_),
    .B(_11737_),
    .C(_11739_),
    .D(_11744_),
    .X(_11745_));
 sky130_fd_sc_hd__nor2_1 _16026_ (.A(_11735_),
    .B(_11745_),
    .Y(_11746_));
 sky130_fd_sc_hd__and2b_1 _16027_ (.A_N(_09987_),
    .B(\line_cache[256][6] ),
    .X(_11747_));
 sky130_fd_sc_hd__and2b_1 _16028_ (.A_N(_09747_),
    .B(\line_cache[302][6] ),
    .X(_11748_));
 sky130_fd_sc_hd__a22o_1 _16029_ (.A1(_09743_),
    .A2(\line_cache[301][6] ),
    .B1(\line_cache[300][6] ),
    .B2(_09742_),
    .X(_11749_));
 sky130_fd_sc_hd__or3_1 _16030_ (.A(_11747_),
    .B(_11748_),
    .C(_11749_),
    .X(_11750_));
 sky130_fd_sc_hd__and3_1 _16031_ (.A(_09917_),
    .B(_09546_),
    .C(\line_cache[258][6] ),
    .X(_11751_));
 sky130_fd_sc_hd__and3_1 _16032_ (.A(_09848_),
    .B(_09691_),
    .C(\line_cache[260][6] ),
    .X(_11752_));
 sky130_fd_sc_hd__and3_1 _16033_ (.A(_09919_),
    .B(_09691_),
    .C(\line_cache[257][6] ),
    .X(_11753_));
 sky130_fd_sc_hd__and3_1 _16034_ (.A(_09840_),
    .B(_09611_),
    .C(\line_cache[259][6] ),
    .X(_11754_));
 sky130_fd_sc_hd__or4_1 _16035_ (.A(_11751_),
    .B(_11752_),
    .C(_11753_),
    .D(_11754_),
    .X(_11755_));
 sky130_fd_sc_hd__and3_1 _16036_ (.A(_09858_),
    .B(_09547_),
    .C(\line_cache[267][6] ),
    .X(_11756_));
 sky130_fd_sc_hd__a22o_1 _16037_ (.A1(_09998_),
    .A2(\line_cache[265][6] ),
    .B1(\line_cache[266][6] ),
    .B2(_09999_),
    .X(_11757_));
 sky130_fd_sc_hd__a311o_1 _16038_ (.A1(_09548_),
    .A2(\line_cache[268][6] ),
    .A3(_09862_),
    .B1(_11756_),
    .C1(_11757_),
    .X(_11758_));
 sky130_fd_sc_hd__nand2_1 _16039_ (.A(_10007_),
    .B(\line_cache[262][6] ),
    .Y(_11759_));
 sky130_fd_sc_hd__nand2_1 _16040_ (.A(_10010_),
    .B(\line_cache[261][6] ),
    .Y(_11760_));
 sky130_fd_sc_hd__nand2_1 _16041_ (.A(_11759_),
    .B(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__a221oi_1 _16042_ (.A1(_10003_),
    .A2(\line_cache[264][6] ),
    .B1(_10005_),
    .B2(\line_cache[263][6] ),
    .C1(_11761_),
    .Y(_11762_));
 sky130_fd_sc_hd__or4b_1 _16043_ (.A(_11750_),
    .B(_11755_),
    .C(_11758_),
    .D_N(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__a22o_1 _16044_ (.A1(_09682_),
    .A2(\line_cache[308][6] ),
    .B1(\line_cache[309][6] ),
    .B2(_09685_),
    .X(_11764_));
 sky130_fd_sc_hd__a221o_1 _16045_ (.A1(\line_cache[311][6] ),
    .A2(_09689_),
    .B1(\line_cache[310][6] ),
    .B2(_09693_),
    .C1(_11764_),
    .X(_11765_));
 sky130_fd_sc_hd__a22o_1 _16046_ (.A1(_09728_),
    .A2(\line_cache[295][6] ),
    .B1(\line_cache[294][6] ),
    .B2(_09726_),
    .X(_11766_));
 sky130_fd_sc_hd__a221o_1 _16047_ (.A1(\line_cache[293][6] ),
    .A2(_09730_),
    .B1(\line_cache[292][6] ),
    .B2(_10018_),
    .C1(_11766_),
    .X(_11767_));
 sky130_fd_sc_hd__a22o_1 _16048_ (.A1(_09716_),
    .A2(\line_cache[296][6] ),
    .B1(\line_cache[297][6] ),
    .B2(_09721_),
    .X(_11768_));
 sky130_fd_sc_hd__a221o_1 _16049_ (.A1(\line_cache[299][6] ),
    .A2(_09718_),
    .B1(\line_cache[298][6] ),
    .B2(_09720_),
    .C1(_11768_),
    .X(_11769_));
 sky130_fd_sc_hd__a22o_1 _16050_ (.A1(_10025_),
    .A2(\line_cache[288][6] ),
    .B1(\line_cache[289][6] ),
    .B2(_10026_),
    .X(_11770_));
 sky130_fd_sc_hd__a221o_1 _16051_ (.A1(\line_cache[291][6] ),
    .A2(_10023_),
    .B1(\line_cache[290][6] ),
    .B2(_10024_),
    .C1(_11770_),
    .X(_11771_));
 sky130_fd_sc_hd__or4_2 _16052_ (.A(_11765_),
    .B(_11767_),
    .C(_11769_),
    .D(_11771_),
    .X(_11772_));
 sky130_fd_sc_hd__nor2_1 _16053_ (.A(_11763_),
    .B(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand2_1 _16054_ (.A(_11746_),
    .B(_11773_),
    .Y(_11774_));
 sky130_fd_sc_hd__nor2_1 _16055_ (.A(_11722_),
    .B(_11774_),
    .Y(_11775_));
 sky130_fd_sc_hd__a22o_1 _16056_ (.A1(_09842_),
    .A2(\line_cache[6][6] ),
    .B1(\line_cache[5][6] ),
    .B2(_09844_),
    .X(_11776_));
 sky130_fd_sc_hd__a221o_1 _16057_ (.A1(\line_cache[4][6] ),
    .A2(_09850_),
    .B1(\line_cache[3][6] ),
    .B2(_09914_),
    .C1(_11776_),
    .X(_11777_));
 sky130_fd_sc_hd__and3_1 _16058_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][6] ),
    .X(_11778_));
 sky130_fd_sc_hd__and3_1 _16059_ (.A(_09919_),
    .B(_09533_),
    .C(\line_cache[1][6] ),
    .X(_11779_));
 sky130_fd_sc_hd__a211o_1 _16060_ (.A1(\line_cache[15][6] ),
    .A2(_09867_),
    .B1(_11778_),
    .C1(_11779_),
    .X(_11780_));
 sky130_fd_sc_hd__and3_1 _16061_ (.A(_09922_),
    .B(_09531_),
    .C(\line_cache[63][6] ),
    .X(_11781_));
 sky130_fd_sc_hd__a31o_1 _16062_ (.A1(_09547_),
    .A2(\line_cache[319][6] ),
    .A3(_09922_),
    .B1(_11781_),
    .X(_11782_));
 sky130_fd_sc_hd__a221o_1 _16063_ (.A1(\line_cache[47][6] ),
    .A2(_09806_),
    .B1(\line_cache[31][6] ),
    .B2(_09907_),
    .C1(_11782_),
    .X(_11783_));
 sky130_fd_sc_hd__nand2_1 _16064_ (.A(_09746_),
    .B(\line_cache[303][6] ),
    .Y(_11784_));
 sky130_fd_sc_hd__nand2_1 _16065_ (.A(_09930_),
    .B(\line_cache[271][6] ),
    .Y(_11785_));
 sky130_fd_sc_hd__nand2_1 _16066_ (.A(_11784_),
    .B(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__a221oi_2 _16067_ (.A1(\line_cache[255][6] ),
    .A2(_09926_),
    .B1(\line_cache[287][6] ),
    .B2(_09927_),
    .C1(_11786_),
    .Y(_11787_));
 sky130_fd_sc_hd__or4b_1 _16068_ (.A(_11777_),
    .B(_11780_),
    .C(_11783_),
    .D_N(_11787_),
    .X(_11788_));
 sky130_fd_sc_hd__a22o_1 _16069_ (.A1(_09803_),
    .A2(\line_cache[45][6] ),
    .B1(\line_cache[46][6] ),
    .B2(_09804_),
    .X(_11789_));
 sky130_fd_sc_hd__a22o_1 _16070_ (.A1(_09824_),
    .A2(\line_cache[48][6] ),
    .B1(\line_cache[49][6] ),
    .B2(_09826_),
    .X(_11790_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_09787_),
    .B(\line_cache[41][6] ),
    .Y(_11791_));
 sky130_fd_sc_hd__nand2_1 _16072_ (.A(_09789_),
    .B(\line_cache[42][6] ),
    .Y(_11792_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(_11791_),
    .B(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__a221oi_2 _16074_ (.A1(_09785_),
    .A2(\line_cache[43][6] ),
    .B1(\line_cache[44][6] ),
    .B2(_09801_),
    .C1(_11793_),
    .Y(_11794_));
 sky130_fd_sc_hd__or3b_1 _16075_ (.A(_11789_),
    .B(_11790_),
    .C_N(_11794_),
    .X(_11795_));
 sky130_fd_sc_hd__a22o_1 _16076_ (.A1(_09699_),
    .A2(\line_cache[317][6] ),
    .B1(\line_cache[316][6] ),
    .B2(_09697_),
    .X(_11796_));
 sky130_fd_sc_hd__a22o_1 _16077_ (.A1(_09832_),
    .A2(\line_cache[58][6] ),
    .B1(\line_cache[59][6] ),
    .B2(_09833_),
    .X(_11797_));
 sky130_fd_sc_hd__a22o_1 _16078_ (.A1(_09819_),
    .A2(\line_cache[61][6] ),
    .B1(\line_cache[60][6] ),
    .B2(_09817_),
    .X(_11798_));
 sky130_fd_sc_hd__a22o_1 _16079_ (.A1(_09822_),
    .A2(\line_cache[62][6] ),
    .B1(\line_cache[318][6] ),
    .B2(_09702_),
    .X(_11799_));
 sky130_fd_sc_hd__or4_1 _16080_ (.A(_11796_),
    .B(_11797_),
    .C(_11798_),
    .D(_11799_),
    .X(_11800_));
 sky130_fd_sc_hd__a22o_1 _16081_ (.A1(_09675_),
    .A2(\line_cache[304][6] ),
    .B1(\line_cache[305][6] ),
    .B2(_09676_),
    .X(_11801_));
 sky130_fd_sc_hd__a22o_1 _16082_ (.A1(_09705_),
    .A2(\line_cache[312][6] ),
    .B1(\line_cache[313][6] ),
    .B2(_09707_),
    .X(_11802_));
 sky130_fd_sc_hd__a22o_1 _16083_ (.A1(_09708_),
    .A2(\line_cache[314][6] ),
    .B1(\line_cache[315][6] ),
    .B2(_09709_),
    .X(_11803_));
 sky130_fd_sc_hd__a22o_1 _16084_ (.A1(_09677_),
    .A2(\line_cache[306][6] ),
    .B1(\line_cache[307][6] ),
    .B2(_09678_),
    .X(_11804_));
 sky130_fd_sc_hd__or4_1 _16085_ (.A(_11801_),
    .B(_11802_),
    .C(_11803_),
    .D(_11804_),
    .X(_11805_));
 sky130_fd_sc_hd__a22o_1 _16086_ (.A1(_09830_),
    .A2(\line_cache[56][6] ),
    .B1(\line_cache[57][6] ),
    .B2(_09834_),
    .X(_11806_));
 sky130_fd_sc_hd__a22o_1 _16087_ (.A1(_09809_),
    .A2(\line_cache[52][6] ),
    .B1(\line_cache[53][6] ),
    .B2(_09811_),
    .X(_11807_));
 sky130_fd_sc_hd__a22o_1 _16088_ (.A1(_09827_),
    .A2(\line_cache[50][6] ),
    .B1(\line_cache[51][6] ),
    .B2(_09828_),
    .X(_11808_));
 sky130_fd_sc_hd__a22o_1 _16089_ (.A1(_09813_),
    .A2(\line_cache[54][6] ),
    .B1(\line_cache[55][6] ),
    .B2(_09815_),
    .X(_11809_));
 sky130_fd_sc_hd__or4_1 _16090_ (.A(_11806_),
    .B(_11807_),
    .C(_11808_),
    .D(_11809_),
    .X(_11810_));
 sky130_fd_sc_hd__or4_2 _16091_ (.A(_11795_),
    .B(_11800_),
    .C(_11805_),
    .D(_11810_),
    .X(_11811_));
 sky130_fd_sc_hd__nand2_1 _16092_ (.A(_09864_),
    .B(\line_cache[12][6] ),
    .Y(_11812_));
 sky130_fd_sc_hd__nand2_1 _16093_ (.A(_09860_),
    .B(\line_cache[11][6] ),
    .Y(_11813_));
 sky130_fd_sc_hd__nand2_1 _16094_ (.A(_11812_),
    .B(_11813_),
    .Y(_11814_));
 sky130_fd_sc_hd__a221oi_2 _16095_ (.A1(_09870_),
    .A2(\line_cache[14][6] ),
    .B1(\line_cache[13][6] ),
    .B2(_09873_),
    .C1(_11814_),
    .Y(_11815_));
 sky130_fd_sc_hd__nand2_1 _16096_ (.A(_09853_),
    .B(\line_cache[10][6] ),
    .Y(_11816_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(_09857_),
    .B(\line_cache[9][6] ),
    .Y(_11817_));
 sky130_fd_sc_hd__nand2_1 _16098_ (.A(_11816_),
    .B(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__a221oi_1 _16099_ (.A1(_09855_),
    .A2(\line_cache[8][6] ),
    .B1(_09847_),
    .B2(\line_cache[7][6] ),
    .C1(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__nand2_1 _16100_ (.A(_11815_),
    .B(_11819_),
    .Y(_11820_));
 sky130_fd_sc_hd__and3_1 _16101_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][6] ),
    .X(_11821_));
 sky130_fd_sc_hd__a22o_1 _16102_ (.A1(_09884_),
    .A2(\line_cache[23][6] ),
    .B1(\line_cache[22][6] ),
    .B2(_09886_),
    .X(_11822_));
 sky130_fd_sc_hd__a22o_1 _16103_ (.A1(_09877_),
    .A2(\line_cache[19][6] ),
    .B1(\line_cache[18][6] ),
    .B2(_09878_),
    .X(_11823_));
 sky130_fd_sc_hd__a221o_1 _16104_ (.A1(\line_cache[17][6] ),
    .A2(_09969_),
    .B1(\line_cache[16][6] ),
    .B2(_09970_),
    .C1(_11823_),
    .X(_11824_));
 sky130_fd_sc_hd__a2111o_1 _16105_ (.A1(\line_cache[20][6] ),
    .A2(_09888_),
    .B1(_11821_),
    .C1(_11822_),
    .D1(_11824_),
    .X(_11825_));
 sky130_fd_sc_hd__a22o_1 _16106_ (.A1(_09796_),
    .A2(\line_cache[33][6] ),
    .B1(\line_cache[34][6] ),
    .B2(_09798_),
    .X(_11826_));
 sky130_fd_sc_hd__a221o_1 _16107_ (.A1(\line_cache[36][6] ),
    .A2(_09777_),
    .B1(\line_cache[35][6] ),
    .B2(_09794_),
    .C1(_11826_),
    .X(_11827_));
 sky130_fd_sc_hd__a22o_1 _16108_ (.A1(_09890_),
    .A2(\line_cache[27][6] ),
    .B1(\line_cache[26][6] ),
    .B2(_09896_),
    .X(_11828_));
 sky130_fd_sc_hd__a221oi_1 _16109_ (.A1(\line_cache[25][6] ),
    .A2(_09892_),
    .B1(\line_cache[24][6] ),
    .B2(_09895_),
    .C1(_11828_),
    .Y(_11829_));
 sky130_fd_sc_hd__a22o_1 _16110_ (.A1(_09903_),
    .A2(\line_cache[29][6] ),
    .B1(\line_cache[28][6] ),
    .B2(_09900_),
    .X(_11830_));
 sky130_fd_sc_hd__a221oi_1 _16111_ (.A1(\line_cache[32][6] ),
    .A2(_09792_),
    .B1(\line_cache[30][6] ),
    .B2(_09905_),
    .C1(_11830_),
    .Y(_11831_));
 sky130_fd_sc_hd__nand2_1 _16112_ (.A(_09773_),
    .B(\line_cache[38][6] ),
    .Y(_11832_));
 sky130_fd_sc_hd__nand2_1 _16113_ (.A(_09775_),
    .B(\line_cache[37][6] ),
    .Y(_11833_));
 sky130_fd_sc_hd__nand2_1 _16114_ (.A(_11832_),
    .B(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__a221oi_4 _16115_ (.A1(_09783_),
    .A2(\line_cache[40][6] ),
    .B1(\line_cache[39][6] ),
    .B2(_09780_),
    .C1(_11834_),
    .Y(_11835_));
 sky130_fd_sc_hd__and4b_1 _16116_ (.A_N(_11827_),
    .B(_11829_),
    .C(_11831_),
    .D(_11835_),
    .X(_11836_));
 sky130_fd_sc_hd__or3b_1 _16117_ (.A(_11820_),
    .B(_11825_),
    .C_N(_11836_),
    .X(_11837_));
 sky130_fd_sc_hd__nor3_2 _16118_ (.A(_11788_),
    .B(_11811_),
    .C(_11837_),
    .Y(_11838_));
 sky130_fd_sc_hd__a22o_1 _16119_ (.A1(_10244_),
    .A2(\line_cache[173][6] ),
    .B1(\line_cache[172][6] ),
    .B2(_10245_),
    .X(_11839_));
 sky130_fd_sc_hd__a221o_1 _16120_ (.A1(\line_cache[175][6] ),
    .A2(_10242_),
    .B1(\line_cache[174][6] ),
    .B2(_10243_),
    .C1(_11839_),
    .X(_11840_));
 sky130_fd_sc_hd__a22o_1 _16121_ (.A1(_10263_),
    .A2(\line_cache[170][6] ),
    .B1(\line_cache[171][6] ),
    .B2(_10262_),
    .X(_11841_));
 sky130_fd_sc_hd__a221o_1 _16122_ (.A1(\line_cache[169][6] ),
    .A2(_10260_),
    .B1(\line_cache[168][6] ),
    .B2(_10261_),
    .C1(_11841_),
    .X(_11842_));
 sky130_fd_sc_hd__a22o_1 _16123_ (.A1(_10256_),
    .A2(\line_cache[160][6] ),
    .B1(\line_cache[161][6] ),
    .B2(_10257_),
    .X(_11843_));
 sky130_fd_sc_hd__and3_1 _16124_ (.A(_10104_),
    .B(_09751_),
    .C(\line_cache[163][6] ),
    .X(_11844_));
 sky130_fd_sc_hd__a22o_1 _16125_ (.A1(_10249_),
    .A2(\line_cache[166][6] ),
    .B1(\line_cache[167][6] ),
    .B2(_10248_),
    .X(_11845_));
 sky130_fd_sc_hd__a221o_1 _16126_ (.A1(\line_cache[165][6] ),
    .A2(_10250_),
    .B1(\line_cache[164][6] ),
    .B2(_10251_),
    .C1(_11845_),
    .X(_11846_));
 sky130_fd_sc_hd__a2111o_1 _16127_ (.A1(\line_cache[162][6] ),
    .A2(_10255_),
    .B1(_11843_),
    .C1(_11844_),
    .D1(_11846_),
    .X(_11847_));
 sky130_fd_sc_hd__nor3_1 _16128_ (.A(_11840_),
    .B(_11842_),
    .C(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__a22o_1 _16129_ (.A1(_10272_),
    .A2(\line_cache[189][6] ),
    .B1(\line_cache[188][6] ),
    .B2(_10271_),
    .X(_11849_));
 sky130_fd_sc_hd__a221o_1 _16130_ (.A1(\line_cache[191][6] ),
    .A2(_10269_),
    .B1(\line_cache[190][6] ),
    .B2(_10270_),
    .C1(_11849_),
    .X(_11850_));
 sky130_fd_sc_hd__a22o_1 _16131_ (.A1(_10284_),
    .A2(\line_cache[176][6] ),
    .B1(_10285_),
    .B2(\line_cache[177][6] ),
    .X(_11851_));
 sky130_fd_sc_hd__a221oi_2 _16132_ (.A1(\line_cache[179][6] ),
    .A2(_10282_),
    .B1(\line_cache[178][6] ),
    .B2(_10283_),
    .C1(_11851_),
    .Y(_11852_));
 sky130_fd_sc_hd__and3_1 _16133_ (.A(_10288_),
    .B(_10102_),
    .C(\line_cache[182][6] ),
    .X(_11853_));
 sky130_fd_sc_hd__and3_1 _16134_ (.A(_10288_),
    .B(_10098_),
    .C(\line_cache[181][6] ),
    .X(_11854_));
 sky130_fd_sc_hd__a31o_1 _16135_ (.A1(\line_cache[180][6] ),
    .A2(_10289_),
    .A3(_10106_),
    .B1(_11854_),
    .X(_11855_));
 sky130_fd_sc_hd__a311oi_2 _16136_ (.A1(\line_cache[183][6] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_11853_),
    .C1(_11855_),
    .Y(_11856_));
 sky130_fd_sc_hd__a22o_1 _16137_ (.A1(_10277_),
    .A2(\line_cache[184][6] ),
    .B1(\line_cache[185][6] ),
    .B2(_10278_),
    .X(_11857_));
 sky130_fd_sc_hd__a221oi_2 _16138_ (.A1(\line_cache[187][6] ),
    .A2(_10275_),
    .B1(\line_cache[186][6] ),
    .B2(_10276_),
    .C1(_11857_),
    .Y(_11858_));
 sky130_fd_sc_hd__and4b_1 _16139_ (.A_N(_11850_),
    .B(_11852_),
    .C(_11856_),
    .D(_11858_),
    .X(_11859_));
 sky130_fd_sc_hd__a22o_1 _16140_ (.A1(_10219_),
    .A2(\line_cache[157][6] ),
    .B1(\line_cache[156][6] ),
    .B2(_10220_),
    .X(_11860_));
 sky130_fd_sc_hd__a221o_1 _16141_ (.A1(\line_cache[159][6] ),
    .A2(_10217_),
    .B1(\line_cache[158][6] ),
    .B2(_10218_),
    .C1(_11860_),
    .X(_11861_));
 sky130_fd_sc_hd__a22o_1 _16142_ (.A1(_10225_),
    .A2(\line_cache[151][6] ),
    .B1(\line_cache[150][6] ),
    .B2(_10226_),
    .X(_11862_));
 sky130_fd_sc_hd__a221oi_2 _16143_ (.A1(\line_cache[149][6] ),
    .A2(_10223_),
    .B1(\line_cache[148][6] ),
    .B2(_10224_),
    .C1(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__a22o_1 _16144_ (.A1(_10231_),
    .A2(\line_cache[147][6] ),
    .B1(\line_cache[146][6] ),
    .B2(_10232_),
    .X(_11864_));
 sky130_fd_sc_hd__a221oi_2 _16145_ (.A1(\line_cache[145][6] ),
    .A2(_10229_),
    .B1(\line_cache[144][6] ),
    .B2(_10230_),
    .C1(_11864_),
    .Y(_11865_));
 sky130_fd_sc_hd__a22o_1 _16146_ (.A1(_10237_),
    .A2(\line_cache[155][6] ),
    .B1(\line_cache[154][6] ),
    .B2(_10238_),
    .X(_11866_));
 sky130_fd_sc_hd__a221oi_1 _16147_ (.A1(\line_cache[153][6] ),
    .A2(_10235_),
    .B1(\line_cache[152][6] ),
    .B2(_10236_),
    .C1(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__and4b_1 _16148_ (.A_N(_11861_),
    .B(_11863_),
    .C(_11865_),
    .D(_11867_),
    .X(_11868_));
 sky130_fd_sc_hd__and3_2 _16149_ (.A(_11848_),
    .B(_11859_),
    .C(_11868_),
    .X(_11869_));
 sky130_fd_sc_hd__a22o_1 _16150_ (.A1(_10378_),
    .A2(\line_cache[80][6] ),
    .B1(_10379_),
    .B2(\line_cache[81][6] ),
    .X(_11870_));
 sky130_fd_sc_hd__a221o_1 _16151_ (.A1(\line_cache[83][6] ),
    .A2(_10376_),
    .B1(\line_cache[82][6] ),
    .B2(_10377_),
    .C1(_11870_),
    .X(_11871_));
 sky130_fd_sc_hd__a22o_1 _16152_ (.A1(_10384_),
    .A2(\line_cache[92][6] ),
    .B1(_10385_),
    .B2(\line_cache[93][6] ),
    .X(_11872_));
 sky130_fd_sc_hd__a221o_1 _16153_ (.A1(\line_cache[95][6] ),
    .A2(net136),
    .B1(\line_cache[94][6] ),
    .B2(_10383_),
    .C1(_11872_),
    .X(_11873_));
 sky130_fd_sc_hd__a22o_1 _16154_ (.A1(_10390_),
    .A2(\line_cache[84][6] ),
    .B1(_10391_),
    .B2(\line_cache[85][6] ),
    .X(_11874_));
 sky130_fd_sc_hd__a221o_1 _16155_ (.A1(\line_cache[87][6] ),
    .A2(_10388_),
    .B1(\line_cache[86][6] ),
    .B2(_10389_),
    .C1(_11874_),
    .X(_11875_));
 sky130_fd_sc_hd__a22o_1 _16156_ (.A1(_10396_),
    .A2(\line_cache[88][6] ),
    .B1(_10397_),
    .B2(\line_cache[89][6] ),
    .X(_11876_));
 sky130_fd_sc_hd__a221o_1 _16157_ (.A1(\line_cache[91][6] ),
    .A2(_10394_),
    .B1(\line_cache[90][6] ),
    .B2(_10395_),
    .C1(_11876_),
    .X(_11877_));
 sky130_fd_sc_hd__or4_1 _16158_ (.A(_11871_),
    .B(_11873_),
    .C(_11875_),
    .D(_11877_),
    .X(_11878_));
 sky130_fd_sc_hd__a22o_1 _16159_ (.A1(_10371_),
    .A2(\line_cache[100][6] ),
    .B1(_10372_),
    .B2(\line_cache[101][6] ),
    .X(_11879_));
 sky130_fd_sc_hd__a22o_1 _16160_ (.A1(_10369_),
    .A2(\line_cache[103][6] ),
    .B1(_10370_),
    .B2(\line_cache[102][6] ),
    .X(_11880_));
 sky130_fd_sc_hd__a22o_1 _16161_ (.A1(_10351_),
    .A2(\line_cache[96][6] ),
    .B1(_10352_),
    .B2(\line_cache[97][6] ),
    .X(_11881_));
 sky130_fd_sc_hd__a221o_2 _16162_ (.A1(\line_cache[99][6] ),
    .A2(_10349_),
    .B1(\line_cache[98][6] ),
    .B2(_10348_),
    .C1(_11881_),
    .X(_11882_));
 sky130_fd_sc_hd__and3_1 _16163_ (.A(_10035_),
    .B(\line_cache[107][6] ),
    .C(_10651_),
    .X(_11883_));
 sky130_fd_sc_hd__and3_1 _16164_ (.A(_10176_),
    .B(\line_cache[105][6] ),
    .C(_10651_),
    .X(_11884_));
 sky130_fd_sc_hd__and3_1 _16165_ (.A(_10054_),
    .B(\line_cache[106][6] ),
    .C(_10356_),
    .X(_11885_));
 sky130_fd_sc_hd__and3_1 _16166_ (.A(_10360_),
    .B(\line_cache[104][6] ),
    .C(_10356_),
    .X(_11886_));
 sky130_fd_sc_hd__or4_1 _16167_ (.A(_11883_),
    .B(_11884_),
    .C(_11885_),
    .D(_11886_),
    .X(_11887_));
 sky130_fd_sc_hd__a22o_1 _16168_ (.A1(_10365_),
    .A2(\line_cache[108][6] ),
    .B1(_10366_),
    .B2(\line_cache[109][6] ),
    .X(_11888_));
 sky130_fd_sc_hd__a221o_1 _16169_ (.A1(\line_cache[111][6] ),
    .A2(_10363_),
    .B1(\line_cache[110][6] ),
    .B2(_10364_),
    .C1(_11888_),
    .X(_11889_));
 sky130_fd_sc_hd__or2_1 _16170_ (.A(_11887_),
    .B(_11889_),
    .X(_11890_));
 sky130_fd_sc_hd__or4_1 _16171_ (.A(_11879_),
    .B(_11880_),
    .C(_11882_),
    .D(_11890_),
    .X(_11891_));
 sky130_fd_sc_hd__nor2_1 _16172_ (.A(_11878_),
    .B(_11891_),
    .Y(_11892_));
 sky130_fd_sc_hd__and3_1 _16173_ (.A(_09758_),
    .B(_10031_),
    .C(\line_cache[141][6] ),
    .X(_11893_));
 sky130_fd_sc_hd__a21o_1 _16174_ (.A1(\line_cache[140][6] ),
    .A2(_10336_),
    .B1(_11893_),
    .X(_11894_));
 sky130_fd_sc_hd__a221o_1 _16175_ (.A1(\line_cache[143][6] ),
    .A2(_10334_),
    .B1(\line_cache[142][6] ),
    .B2(_10335_),
    .C1(_11894_),
    .X(_11895_));
 sky130_fd_sc_hd__and3_1 _16176_ (.A(_09758_),
    .B(_10098_),
    .C(\line_cache[133][6] ),
    .X(_11896_));
 sky130_fd_sc_hd__a21o_1 _16177_ (.A1(\line_cache[132][6] ),
    .A2(_10324_),
    .B1(_11896_),
    .X(_11897_));
 sky130_fd_sc_hd__a221o_1 _16178_ (.A1(\line_cache[135][6] ),
    .A2(_10322_),
    .B1(\line_cache[134][6] ),
    .B2(_10323_),
    .C1(_11897_),
    .X(_11898_));
 sky130_fd_sc_hd__and3_1 _16179_ (.A(_10071_),
    .B(\line_cache[128][6] ),
    .C(_09758_),
    .X(_11899_));
 sky130_fd_sc_hd__a21o_1 _16180_ (.A1(\line_cache[129][6] ),
    .A2(_10330_),
    .B1(_11899_),
    .X(_11900_));
 sky130_fd_sc_hd__a221o_1 _16181_ (.A1(\line_cache[131][6] ),
    .A2(_10328_),
    .B1(\line_cache[130][6] ),
    .B2(_10329_),
    .C1(_11900_),
    .X(_11901_));
 sky130_fd_sc_hd__a22o_1 _16182_ (.A1(_10342_),
    .A2(\line_cache[139][6] ),
    .B1(\line_cache[138][6] ),
    .B2(_10343_),
    .X(_11902_));
 sky130_fd_sc_hd__a221o_1 _16183_ (.A1(\line_cache[137][6] ),
    .A2(_10340_),
    .B1(\line_cache[136][6] ),
    .B2(_10341_),
    .C1(_11902_),
    .X(_11903_));
 sky130_fd_sc_hd__or4_1 _16184_ (.A(_11895_),
    .B(_11898_),
    .C(_11901_),
    .D(_11903_),
    .X(_11904_));
 sky130_fd_sc_hd__a22o_1 _16185_ (.A1(_10298_),
    .A2(\line_cache[112][6] ),
    .B1(_10299_),
    .B2(\line_cache[113][6] ),
    .X(_11905_));
 sky130_fd_sc_hd__a221o_1 _16186_ (.A1(\line_cache[115][6] ),
    .A2(_10296_),
    .B1(\line_cache[114][6] ),
    .B2(_10297_),
    .C1(_11905_),
    .X(_11906_));
 sky130_fd_sc_hd__a22o_1 _16187_ (.A1(_10305_),
    .A2(\line_cache[124][6] ),
    .B1(_10306_),
    .B2(\line_cache[125][6] ),
    .X(_11907_));
 sky130_fd_sc_hd__a221o_1 _16188_ (.A1(\line_cache[126][6] ),
    .A2(_10304_),
    .B1(\line_cache[127][6] ),
    .B2(_10622_),
    .C1(_11907_),
    .X(_11908_));
 sky130_fd_sc_hd__a22o_1 _16189_ (.A1(_10311_),
    .A2(\line_cache[116][6] ),
    .B1(_10312_),
    .B2(\line_cache[117][6] ),
    .X(_11909_));
 sky130_fd_sc_hd__a221o_1 _16190_ (.A1(\line_cache[119][6] ),
    .A2(_10309_),
    .B1(\line_cache[118][6] ),
    .B2(_10310_),
    .C1(_11909_),
    .X(_11910_));
 sky130_fd_sc_hd__a22o_1 _16191_ (.A1(_10317_),
    .A2(\line_cache[120][6] ),
    .B1(_10318_),
    .B2(\line_cache[121][6] ),
    .X(_11911_));
 sky130_fd_sc_hd__a221o_1 _16192_ (.A1(\line_cache[123][6] ),
    .A2(_10315_),
    .B1(\line_cache[122][6] ),
    .B2(_10316_),
    .C1(_11911_),
    .X(_11912_));
 sky130_fd_sc_hd__or4_1 _16193_ (.A(_11906_),
    .B(_11908_),
    .C(_11910_),
    .D(_11912_),
    .X(_11913_));
 sky130_fd_sc_hd__nor2_1 _16194_ (.A(_11904_),
    .B(_11913_),
    .Y(_11914_));
 sky130_fd_sc_hd__and3_1 _16195_ (.A(_11869_),
    .B(_11892_),
    .C(_11914_),
    .X(_11915_));
 sky130_fd_sc_hd__nand3_1 _16196_ (.A(_11775_),
    .B(_11838_),
    .C(_11915_),
    .Y(_11916_));
 sky130_fd_sc_hd__o21ba_2 _16197_ (.A1(_11668_),
    .A2(_11916_),
    .B1_N(_08979_),
    .X(_11917_));
 sky130_fd_sc_hd__buf_6 _16198_ (.A(_11917_),
    .X(net132));
 sky130_fd_sc_hd__and2_1 _16199_ (.A(_09912_),
    .B(\line_cache[0][7] ),
    .X(_11918_));
 sky130_fd_sc_hd__and3_1 _16200_ (.A(_10031_),
    .B(\line_cache[77][7] ),
    .C(_10167_),
    .X(_11919_));
 sky130_fd_sc_hd__and3_1 _16201_ (.A(_10038_),
    .B(\line_cache[78][7] ),
    .C(_10167_),
    .X(_11920_));
 sky130_fd_sc_hd__and3_1 _16202_ (.A(_10041_),
    .B(\line_cache[76][7] ),
    .C(_10161_),
    .X(_11921_));
 sky130_fd_sc_hd__a2111o_1 _16203_ (.A1(_10168_),
    .A2(\line_cache[79][7] ),
    .B1(_11919_),
    .C1(_11920_),
    .D1(_11921_),
    .X(_11922_));
 sky130_fd_sc_hd__a22o_1 _16204_ (.A1(_10182_),
    .A2(\line_cache[64][7] ),
    .B1(_10183_),
    .B2(\line_cache[65][7] ),
    .X(_11923_));
 sky130_fd_sc_hd__a221o_1 _16205_ (.A1(\line_cache[67][7] ),
    .A2(_10180_),
    .B1(\line_cache[66][7] ),
    .B2(_10181_),
    .C1(_11923_),
    .X(_11924_));
 sky130_fd_sc_hd__a22o_1 _16206_ (.A1(_10163_),
    .A2(\line_cache[68][7] ),
    .B1(_10164_),
    .B2(\line_cache[69][7] ),
    .X(_11925_));
 sky130_fd_sc_hd__a221o_1 _16207_ (.A1(\line_cache[71][7] ),
    .A2(_10159_),
    .B1(\line_cache[70][7] ),
    .B2(_10750_),
    .C1(_11925_),
    .X(_11926_));
 sky130_fd_sc_hd__a22o_1 _16208_ (.A1(_10175_),
    .A2(\line_cache[72][7] ),
    .B1(_10753_),
    .B2(\line_cache[73][7] ),
    .X(_11927_));
 sky130_fd_sc_hd__a221o_1 _16209_ (.A1(\line_cache[75][7] ),
    .A2(_10173_),
    .B1(\line_cache[74][7] ),
    .B2(_10174_),
    .C1(_11927_),
    .X(_11928_));
 sky130_fd_sc_hd__or4_2 _16210_ (.A(_11922_),
    .B(_11924_),
    .C(_11926_),
    .D(_11928_),
    .X(_11929_));
 sky130_fd_sc_hd__a22o_1 _16211_ (.A1(_10189_),
    .A2(\line_cache[252][7] ),
    .B1(_10190_),
    .B2(\line_cache[251][7] ),
    .X(_11930_));
 sky130_fd_sc_hd__a221o_1 _16212_ (.A1(\line_cache[254][7] ),
    .A2(_10187_),
    .B1(\line_cache[253][7] ),
    .B2(_10188_),
    .C1(_11930_),
    .X(_11931_));
 sky130_fd_sc_hd__a22o_1 _16213_ (.A1(_10195_),
    .A2(\line_cache[248][7] ),
    .B1(_10196_),
    .B2(\line_cache[247][7] ),
    .X(_11932_));
 sky130_fd_sc_hd__a221o_1 _16214_ (.A1(\line_cache[250][7] ),
    .A2(_10193_),
    .B1(\line_cache[249][7] ),
    .B2(_10194_),
    .C1(_11932_),
    .X(_11933_));
 sky130_fd_sc_hd__and2b_1 _16215_ (.A_N(_10200_),
    .B(\line_cache[240][7] ),
    .X(_11934_));
 sky130_fd_sc_hd__and2b_1 _16216_ (.A_N(_09570_),
    .B(\line_cache[241][7] ),
    .X(_11935_));
 sky130_fd_sc_hd__and2b_1 _16217_ (.A_N(_10203_),
    .B(\line_cache[242][7] ),
    .X(_11936_));
 sky130_fd_sc_hd__a2111o_1 _16218_ (.A1(\line_cache[239][7] ),
    .A2(_10199_),
    .B1(_11934_),
    .C1(_11935_),
    .D1(_11936_),
    .X(_11937_));
 sky130_fd_sc_hd__and2b_1 _16219_ (.A_N(_10206_),
    .B(\line_cache[243][7] ),
    .X(_11938_));
 sky130_fd_sc_hd__and2b_1 _16220_ (.A_N(_10208_),
    .B(\line_cache[244][7] ),
    .X(_11939_));
 sky130_fd_sc_hd__and2b_1 _16221_ (.A_N(_09597_),
    .B(\line_cache[245][7] ),
    .X(_11940_));
 sky130_fd_sc_hd__and2b_1 _16222_ (.A_N(_10211_),
    .B(\line_cache[246][7] ),
    .X(_11941_));
 sky130_fd_sc_hd__or4_1 _16223_ (.A(_11938_),
    .B(_11939_),
    .C(_11940_),
    .D(_11941_),
    .X(_11942_));
 sky130_fd_sc_hd__or4_1 _16224_ (.A(_11931_),
    .B(_11933_),
    .C(_11937_),
    .D(_11942_),
    .X(_11943_));
 sky130_fd_sc_hd__and3_1 _16225_ (.A(_09595_),
    .B(\line_cache[229][7] ),
    .C(_10099_),
    .X(_11944_));
 sky130_fd_sc_hd__and3_1 _16226_ (.A(_10044_),
    .B(\line_cache[230][7] ),
    .C(_10099_),
    .X(_11945_));
 sky130_fd_sc_hd__and3_1 _16227_ (.A(_10104_),
    .B(\line_cache[227][7] ),
    .C(_10434_),
    .X(_11946_));
 sky130_fd_sc_hd__and3_1 _16228_ (.A(_10106_),
    .B(\line_cache[228][7] ),
    .C(_10437_),
    .X(_11947_));
 sky130_fd_sc_hd__or4_1 _16229_ (.A(_11944_),
    .B(_11945_),
    .C(_11946_),
    .D(_11947_),
    .X(_11948_));
 sky130_fd_sc_hd__and3_1 _16230_ (.A(_09544_),
    .B(\line_cache[223][7] ),
    .C(_09600_),
    .X(_11949_));
 sky130_fd_sc_hd__and3_1 _16231_ (.A(_10070_),
    .B(\line_cache[224][7] ),
    .C(_10434_),
    .X(_11950_));
 sky130_fd_sc_hd__and3_1 _16232_ (.A(_10067_),
    .B(\line_cache[225][7] ),
    .C(_10434_),
    .X(_11951_));
 sky130_fd_sc_hd__and3_1 _16233_ (.A(_10074_),
    .B(\line_cache[226][7] ),
    .C(_10437_),
    .X(_11952_));
 sky130_fd_sc_hd__or4_1 _16234_ (.A(_11949_),
    .B(_11950_),
    .C(_11951_),
    .D(_11952_),
    .X(_11953_));
 sky130_fd_sc_hd__a22o_1 _16235_ (.A1(_10118_),
    .A2(\line_cache[236][7] ),
    .B1(_10120_),
    .B2(\line_cache[235][7] ),
    .X(_11954_));
 sky130_fd_sc_hd__a221o_1 _16236_ (.A1(\line_cache[238][7] ),
    .A2(_10116_),
    .B1(\line_cache[237][7] ),
    .B2(_10117_),
    .C1(_11954_),
    .X(_11955_));
 sky130_fd_sc_hd__a22o_1 _16237_ (.A1(_10125_),
    .A2(\line_cache[232][7] ),
    .B1(_10126_),
    .B2(\line_cache[231][7] ),
    .X(_11956_));
 sky130_fd_sc_hd__a221o_1 _16238_ (.A1(\line_cache[234][7] ),
    .A2(_10123_),
    .B1(\line_cache[233][7] ),
    .B2(_10124_),
    .C1(_11956_),
    .X(_11957_));
 sky130_fd_sc_hd__or4_1 _16239_ (.A(_11948_),
    .B(_11953_),
    .C(_11955_),
    .D(_11957_),
    .X(_11958_));
 sky130_fd_sc_hd__a22o_1 _16240_ (.A1(_10132_),
    .A2(\line_cache[220][7] ),
    .B1(_10133_),
    .B2(\line_cache[219][7] ),
    .X(_11959_));
 sky130_fd_sc_hd__a221o_1 _16241_ (.A1(\line_cache[222][7] ),
    .A2(_10130_),
    .B1(\line_cache[221][7] ),
    .B2(_10131_),
    .C1(_11959_),
    .X(_11960_));
 sky130_fd_sc_hd__a22o_1 _16242_ (.A1(_10138_),
    .A2(\line_cache[208][7] ),
    .B1(_10139_),
    .B2(\line_cache[207][7] ),
    .X(_11961_));
 sky130_fd_sc_hd__a221o_1 _16243_ (.A1(\line_cache[210][7] ),
    .A2(_10136_),
    .B1(\line_cache[209][7] ),
    .B2(_10137_),
    .C1(_11961_),
    .X(_11962_));
 sky130_fd_sc_hd__a22o_1 _16244_ (.A1(_10144_),
    .A2(\line_cache[216][7] ),
    .B1(_10145_),
    .B2(\line_cache[215][7] ),
    .X(_11963_));
 sky130_fd_sc_hd__a221o_1 _16245_ (.A1(\line_cache[218][7] ),
    .A2(_10142_),
    .B1(\line_cache[217][7] ),
    .B2(_10143_),
    .C1(_11963_),
    .X(_11964_));
 sky130_fd_sc_hd__and2b_1 _16246_ (.A_N(_10148_),
    .B(\line_cache[211][7] ),
    .X(_11965_));
 sky130_fd_sc_hd__nor2b_1 _16247_ (.A(_10150_),
    .B_N(\line_cache[212][7] ),
    .Y(_11966_));
 sky130_fd_sc_hd__and2b_1 _16248_ (.A_N(_10152_),
    .B(\line_cache[213][7] ),
    .X(_11967_));
 sky130_fd_sc_hd__and2b_1 _16249_ (.A_N(_10154_),
    .B(\line_cache[214][7] ),
    .X(_11968_));
 sky130_fd_sc_hd__or4_1 _16250_ (.A(_11965_),
    .B(_11966_),
    .C(_11967_),
    .D(_11968_),
    .X(_11969_));
 sky130_fd_sc_hd__or4_2 _16251_ (.A(_11960_),
    .B(_11962_),
    .C(_11964_),
    .D(_11969_),
    .X(_11970_));
 sky130_fd_sc_hd__or2_1 _16252_ (.A(_11958_),
    .B(_11970_),
    .X(_11971_));
 sky130_fd_sc_hd__or3_1 _16253_ (.A(_11929_),
    .B(_11943_),
    .C(_11971_),
    .X(_11972_));
 sky130_fd_sc_hd__and3_1 _16254_ (.A(_10035_),
    .B(\line_cache[203][7] ),
    .C(_09539_),
    .X(_11973_));
 sky130_fd_sc_hd__and3_1 _16255_ (.A(_10038_),
    .B(\line_cache[206][7] ),
    .C(_10075_),
    .X(_11974_));
 sky130_fd_sc_hd__and3_1 _16256_ (.A(_10041_),
    .B(\line_cache[204][7] ),
    .C(_10075_),
    .X(_11975_));
 sky130_fd_sc_hd__a2111o_1 _16257_ (.A1(\line_cache[205][7] ),
    .A2(_10033_),
    .B1(_11973_),
    .C1(_11974_),
    .D1(_11975_),
    .X(_11976_));
 sky130_fd_sc_hd__a22o_1 _16258_ (.A1(_10049_),
    .A2(\line_cache[195][7] ),
    .B1(\line_cache[196][7] ),
    .B2(_10051_),
    .X(_11977_));
 sky130_fd_sc_hd__a221o_1 _16259_ (.A1(\line_cache[198][7] ),
    .A2(_10046_),
    .B1(\line_cache[197][7] ),
    .B2(_10047_),
    .C1(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__a22o_1 _16260_ (.A1(_10060_),
    .A2(\line_cache[200][7] ),
    .B1(_10063_),
    .B2(\line_cache[199][7] ),
    .X(_11979_));
 sky130_fd_sc_hd__a221o_1 _16261_ (.A1(\line_cache[202][7] ),
    .A2(_10056_),
    .B1(\line_cache[201][7] ),
    .B2(_10059_),
    .C1(_11979_),
    .X(_11980_));
 sky130_fd_sc_hd__and3_1 _16262_ (.A(_10067_),
    .B(\line_cache[193][7] ),
    .C(_10075_),
    .X(_11981_));
 sky130_fd_sc_hd__and3_1 _16263_ (.A(_10071_),
    .B(\line_cache[192][7] ),
    .C(_09540_),
    .X(_11982_));
 sky130_fd_sc_hd__and3_1 _16264_ (.A(_10074_),
    .B(\line_cache[194][7] ),
    .C(_09540_),
    .X(_11983_));
 sky130_fd_sc_hd__a2111o_1 _16265_ (.A1(_10066_),
    .A2(\line_cache[286][7] ),
    .B1(_11981_),
    .C1(_11982_),
    .D1(_11983_),
    .X(_11984_));
 sky130_fd_sc_hd__or4_1 _16266_ (.A(_11976_),
    .B(_11978_),
    .C(_11980_),
    .D(_11984_),
    .X(_11985_));
 sky130_fd_sc_hd__a22o_1 _16267_ (.A1(_09623_),
    .A2(\line_cache[275][7] ),
    .B1(_09620_),
    .B2(\line_cache[274][7] ),
    .X(_11986_));
 sky130_fd_sc_hd__a22o_1 _16268_ (.A1(_10080_),
    .A2(\line_cache[276][7] ),
    .B1(\line_cache[277][7] ),
    .B2(_10081_),
    .X(_11987_));
 sky130_fd_sc_hd__a22o_1 _16269_ (.A1(_10086_),
    .A2(\line_cache[270][7] ),
    .B1(\line_cache[269][7] ),
    .B2(_10088_),
    .X(_11988_));
 sky130_fd_sc_hd__a221o_1 _16270_ (.A1(\line_cache[273][7] ),
    .A2(_10083_),
    .B1(\line_cache[272][7] ),
    .B2(_10084_),
    .C1(_11988_),
    .X(_11989_));
 sky130_fd_sc_hd__a22o_1 _16271_ (.A1(_09658_),
    .A2(\line_cache[283][7] ),
    .B1(\line_cache[282][7] ),
    .B2(_09661_),
    .X(_11990_));
 sky130_fd_sc_hd__a22o_1 _16272_ (.A1(_09645_),
    .A2(\line_cache[285][7] ),
    .B1(\line_cache[284][7] ),
    .B2(_09648_),
    .X(_11991_));
 sky130_fd_sc_hd__a22o_1 _16273_ (.A1(_09639_),
    .A2(\line_cache[279][7] ),
    .B1(\line_cache[278][7] ),
    .B2(_09636_),
    .X(_11992_));
 sky130_fd_sc_hd__a221o_1 _16274_ (.A1(\line_cache[281][7] ),
    .A2(_09663_),
    .B1(\line_cache[280][7] ),
    .B2(_09655_),
    .C1(_11992_),
    .X(_11993_));
 sky130_fd_sc_hd__or3_1 _16275_ (.A(_11990_),
    .B(_11991_),
    .C(_11993_),
    .X(_11994_));
 sky130_fd_sc_hd__or4_1 _16276_ (.A(_11986_),
    .B(_11987_),
    .C(_11989_),
    .D(_11994_),
    .X(_11995_));
 sky130_fd_sc_hd__nor2_1 _16277_ (.A(_11985_),
    .B(_11995_),
    .Y(_11996_));
 sky130_fd_sc_hd__and2b_1 _16278_ (.A_N(_09987_),
    .B(\line_cache[256][7] ),
    .X(_11997_));
 sky130_fd_sc_hd__and2b_1 _16279_ (.A_N(_09747_),
    .B(\line_cache[302][7] ),
    .X(_11998_));
 sky130_fd_sc_hd__a22o_1 _16280_ (.A1(_09743_),
    .A2(\line_cache[301][7] ),
    .B1(\line_cache[300][7] ),
    .B2(_09742_),
    .X(_11999_));
 sky130_fd_sc_hd__or3_1 _16281_ (.A(_11997_),
    .B(_11998_),
    .C(_11999_),
    .X(_12000_));
 sky130_fd_sc_hd__and3_1 _16282_ (.A(_09917_),
    .B(_09546_),
    .C(\line_cache[258][7] ),
    .X(_12001_));
 sky130_fd_sc_hd__and3_1 _16283_ (.A(_09848_),
    .B(_09691_),
    .C(\line_cache[260][7] ),
    .X(_12002_));
 sky130_fd_sc_hd__and3_1 _16284_ (.A(_09919_),
    .B(_09691_),
    .C(\line_cache[257][7] ),
    .X(_12003_));
 sky130_fd_sc_hd__and3_1 _16285_ (.A(_09840_),
    .B(_09611_),
    .C(\line_cache[259][7] ),
    .X(_12004_));
 sky130_fd_sc_hd__or4_1 _16286_ (.A(_12001_),
    .B(_12002_),
    .C(_12003_),
    .D(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__and3_1 _16287_ (.A(_09858_),
    .B(_09547_),
    .C(\line_cache[267][7] ),
    .X(_12006_));
 sky130_fd_sc_hd__a22o_1 _16288_ (.A1(_09998_),
    .A2(\line_cache[265][7] ),
    .B1(\line_cache[266][7] ),
    .B2(_09999_),
    .X(_12007_));
 sky130_fd_sc_hd__a311o_1 _16289_ (.A1(_09548_),
    .A2(\line_cache[268][7] ),
    .A3(_09862_),
    .B1(_12006_),
    .C1(_12007_),
    .X(_12008_));
 sky130_fd_sc_hd__nand2_1 _16290_ (.A(_10007_),
    .B(\line_cache[262][7] ),
    .Y(_12009_));
 sky130_fd_sc_hd__nand2_1 _16291_ (.A(_10010_),
    .B(\line_cache[261][7] ),
    .Y(_12010_));
 sky130_fd_sc_hd__nand2_1 _16292_ (.A(_12009_),
    .B(_12010_),
    .Y(_12011_));
 sky130_fd_sc_hd__a221oi_1 _16293_ (.A1(_10003_),
    .A2(\line_cache[264][7] ),
    .B1(_10005_),
    .B2(\line_cache[263][7] ),
    .C1(_12011_),
    .Y(_12012_));
 sky130_fd_sc_hd__or4b_2 _16294_ (.A(_12000_),
    .B(_12005_),
    .C(_12008_),
    .D_N(_12012_),
    .X(_12013_));
 sky130_fd_sc_hd__a22o_1 _16295_ (.A1(_09682_),
    .A2(\line_cache[308][7] ),
    .B1(\line_cache[309][7] ),
    .B2(_09685_),
    .X(_12014_));
 sky130_fd_sc_hd__a221o_1 _16296_ (.A1(\line_cache[311][7] ),
    .A2(_09689_),
    .B1(\line_cache[310][7] ),
    .B2(_09693_),
    .C1(_12014_),
    .X(_12015_));
 sky130_fd_sc_hd__a22o_1 _16297_ (.A1(_09728_),
    .A2(\line_cache[295][7] ),
    .B1(\line_cache[294][7] ),
    .B2(_09726_),
    .X(_12016_));
 sky130_fd_sc_hd__a221o_1 _16298_ (.A1(\line_cache[293][7] ),
    .A2(_09730_),
    .B1(\line_cache[292][7] ),
    .B2(_10018_),
    .C1(_12016_),
    .X(_12017_));
 sky130_fd_sc_hd__a22o_1 _16299_ (.A1(_09716_),
    .A2(\line_cache[296][7] ),
    .B1(\line_cache[297][7] ),
    .B2(_09721_),
    .X(_12018_));
 sky130_fd_sc_hd__a221o_1 _16300_ (.A1(\line_cache[299][7] ),
    .A2(_09718_),
    .B1(\line_cache[298][7] ),
    .B2(_09720_),
    .C1(_12018_),
    .X(_12019_));
 sky130_fd_sc_hd__a22o_1 _16301_ (.A1(_10025_),
    .A2(\line_cache[288][7] ),
    .B1(\line_cache[289][7] ),
    .B2(_10026_),
    .X(_12020_));
 sky130_fd_sc_hd__a221o_1 _16302_ (.A1(\line_cache[291][7] ),
    .A2(_10023_),
    .B1(\line_cache[290][7] ),
    .B2(_10024_),
    .C1(_12020_),
    .X(_12021_));
 sky130_fd_sc_hd__or4_2 _16303_ (.A(_12015_),
    .B(_12017_),
    .C(_12019_),
    .D(_12021_),
    .X(_12022_));
 sky130_fd_sc_hd__nor2_1 _16304_ (.A(_12013_),
    .B(_12022_),
    .Y(_12023_));
 sky130_fd_sc_hd__nand2_1 _16305_ (.A(_11996_),
    .B(_12023_),
    .Y(_12024_));
 sky130_fd_sc_hd__nor2_1 _16306_ (.A(_11972_),
    .B(_12024_),
    .Y(_12025_));
 sky130_fd_sc_hd__a22o_1 _16307_ (.A1(_09842_),
    .A2(\line_cache[6][7] ),
    .B1(\line_cache[5][7] ),
    .B2(_09844_),
    .X(_12026_));
 sky130_fd_sc_hd__a221o_1 _16308_ (.A1(\line_cache[4][7] ),
    .A2(_09850_),
    .B1(\line_cache[3][7] ),
    .B2(_09914_),
    .C1(_12026_),
    .X(_12027_));
 sky130_fd_sc_hd__and3_1 _16309_ (.A(_09917_),
    .B(_09532_),
    .C(\line_cache[2][7] ),
    .X(_12028_));
 sky130_fd_sc_hd__and3_1 _16310_ (.A(_09919_),
    .B(_09532_),
    .C(\line_cache[1][7] ),
    .X(_12029_));
 sky130_fd_sc_hd__a211o_1 _16311_ (.A1(\line_cache[15][7] ),
    .A2(_09867_),
    .B1(_12028_),
    .C1(_12029_),
    .X(_12030_));
 sky130_fd_sc_hd__and3_1 _16312_ (.A(_09922_),
    .B(_09531_),
    .C(\line_cache[63][7] ),
    .X(_12031_));
 sky130_fd_sc_hd__a31o_1 _16313_ (.A1(_09547_),
    .A2(\line_cache[319][7] ),
    .A3(_09922_),
    .B1(_12031_),
    .X(_12032_));
 sky130_fd_sc_hd__a221o_1 _16314_ (.A1(\line_cache[47][7] ),
    .A2(_09806_),
    .B1(\line_cache[31][7] ),
    .B2(_09907_),
    .C1(_12032_),
    .X(_12033_));
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(_09746_),
    .B(\line_cache[303][7] ),
    .Y(_12034_));
 sky130_fd_sc_hd__nand2_1 _16316_ (.A(_09930_),
    .B(\line_cache[271][7] ),
    .Y(_12035_));
 sky130_fd_sc_hd__nand2_1 _16317_ (.A(_12034_),
    .B(_12035_),
    .Y(_12036_));
 sky130_fd_sc_hd__a221oi_2 _16318_ (.A1(\line_cache[255][7] ),
    .A2(_09926_),
    .B1(\line_cache[287][7] ),
    .B2(_09927_),
    .C1(_12036_),
    .Y(_12037_));
 sky130_fd_sc_hd__or4b_1 _16319_ (.A(_12027_),
    .B(_12030_),
    .C(_12033_),
    .D_N(_12037_),
    .X(_12038_));
 sky130_fd_sc_hd__a22o_1 _16320_ (.A1(_09803_),
    .A2(\line_cache[45][7] ),
    .B1(\line_cache[46][7] ),
    .B2(_09804_),
    .X(_12039_));
 sky130_fd_sc_hd__a22o_1 _16321_ (.A1(_09824_),
    .A2(\line_cache[48][7] ),
    .B1(\line_cache[49][7] ),
    .B2(_09826_),
    .X(_12040_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(_09787_),
    .B(\line_cache[41][7] ),
    .Y(_12041_));
 sky130_fd_sc_hd__nand2_1 _16323_ (.A(_09789_),
    .B(\line_cache[42][7] ),
    .Y(_12042_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(_12041_),
    .B(_12042_),
    .Y(_12043_));
 sky130_fd_sc_hd__a221oi_2 _16325_ (.A1(_09785_),
    .A2(\line_cache[43][7] ),
    .B1(\line_cache[44][7] ),
    .B2(_09801_),
    .C1(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__or3b_1 _16326_ (.A(_12039_),
    .B(_12040_),
    .C_N(_12044_),
    .X(_12045_));
 sky130_fd_sc_hd__a22o_1 _16327_ (.A1(_09699_),
    .A2(\line_cache[317][7] ),
    .B1(\line_cache[316][7] ),
    .B2(_09697_),
    .X(_12046_));
 sky130_fd_sc_hd__a22o_1 _16328_ (.A1(_09832_),
    .A2(\line_cache[58][7] ),
    .B1(\line_cache[59][7] ),
    .B2(_09833_),
    .X(_12047_));
 sky130_fd_sc_hd__a22o_1 _16329_ (.A1(_09819_),
    .A2(\line_cache[61][7] ),
    .B1(\line_cache[60][7] ),
    .B2(_09817_),
    .X(_12048_));
 sky130_fd_sc_hd__a22o_1 _16330_ (.A1(_09822_),
    .A2(\line_cache[62][7] ),
    .B1(\line_cache[318][7] ),
    .B2(_09702_),
    .X(_12049_));
 sky130_fd_sc_hd__or4_1 _16331_ (.A(_12046_),
    .B(_12047_),
    .C(_12048_),
    .D(_12049_),
    .X(_12050_));
 sky130_fd_sc_hd__a22o_1 _16332_ (.A1(_09675_),
    .A2(\line_cache[304][7] ),
    .B1(\line_cache[305][7] ),
    .B2(_09676_),
    .X(_12051_));
 sky130_fd_sc_hd__a22o_1 _16333_ (.A1(_09705_),
    .A2(\line_cache[312][7] ),
    .B1(\line_cache[313][7] ),
    .B2(_09707_),
    .X(_12052_));
 sky130_fd_sc_hd__a22o_1 _16334_ (.A1(_09708_),
    .A2(\line_cache[314][7] ),
    .B1(\line_cache[315][7] ),
    .B2(_09709_),
    .X(_12053_));
 sky130_fd_sc_hd__a22o_1 _16335_ (.A1(_09677_),
    .A2(\line_cache[306][7] ),
    .B1(\line_cache[307][7] ),
    .B2(_09678_),
    .X(_12054_));
 sky130_fd_sc_hd__or4_1 _16336_ (.A(_12051_),
    .B(_12052_),
    .C(_12053_),
    .D(_12054_),
    .X(_12055_));
 sky130_fd_sc_hd__a22o_1 _16337_ (.A1(_09830_),
    .A2(\line_cache[56][7] ),
    .B1(\line_cache[57][7] ),
    .B2(_09834_),
    .X(_12056_));
 sky130_fd_sc_hd__a22o_1 _16338_ (.A1(_09809_),
    .A2(\line_cache[52][7] ),
    .B1(\line_cache[53][7] ),
    .B2(_09811_),
    .X(_12057_));
 sky130_fd_sc_hd__a22o_1 _16339_ (.A1(_09827_),
    .A2(\line_cache[50][7] ),
    .B1(\line_cache[51][7] ),
    .B2(_09828_),
    .X(_12058_));
 sky130_fd_sc_hd__a22o_1 _16340_ (.A1(_09813_),
    .A2(\line_cache[54][7] ),
    .B1(\line_cache[55][7] ),
    .B2(_09815_),
    .X(_12059_));
 sky130_fd_sc_hd__or4_1 _16341_ (.A(_12056_),
    .B(_12057_),
    .C(_12058_),
    .D(_12059_),
    .X(_12060_));
 sky130_fd_sc_hd__or4_2 _16342_ (.A(_12045_),
    .B(_12050_),
    .C(_12055_),
    .D(_12060_),
    .X(_12061_));
 sky130_fd_sc_hd__nand2_1 _16343_ (.A(_09864_),
    .B(\line_cache[12][7] ),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_1 _16344_ (.A(_09860_),
    .B(\line_cache[11][7] ),
    .Y(_12063_));
 sky130_fd_sc_hd__nand2_1 _16345_ (.A(_12062_),
    .B(_12063_),
    .Y(_12064_));
 sky130_fd_sc_hd__a221oi_2 _16346_ (.A1(_09870_),
    .A2(\line_cache[14][7] ),
    .B1(\line_cache[13][7] ),
    .B2(_09873_),
    .C1(_12064_),
    .Y(_12065_));
 sky130_fd_sc_hd__nand2_1 _16347_ (.A(_09853_),
    .B(\line_cache[10][7] ),
    .Y(_12066_));
 sky130_fd_sc_hd__nand2_1 _16348_ (.A(_09857_),
    .B(\line_cache[9][7] ),
    .Y(_12067_));
 sky130_fd_sc_hd__nand2_1 _16349_ (.A(_12066_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__a221oi_1 _16350_ (.A1(_09855_),
    .A2(\line_cache[8][7] ),
    .B1(_09847_),
    .B2(\line_cache[7][7] ),
    .C1(_12068_),
    .Y(_12069_));
 sky130_fd_sc_hd__nand2_1 _16351_ (.A(_12065_),
    .B(_12069_),
    .Y(_12070_));
 sky130_fd_sc_hd__and3_1 _16352_ (.A(_09631_),
    .B(_09533_),
    .C(\line_cache[21][7] ),
    .X(_12071_));
 sky130_fd_sc_hd__a22o_1 _16353_ (.A1(_09884_),
    .A2(\line_cache[23][7] ),
    .B1(\line_cache[22][7] ),
    .B2(_09886_),
    .X(_12072_));
 sky130_fd_sc_hd__a22o_1 _16354_ (.A1(_09877_),
    .A2(\line_cache[19][7] ),
    .B1(\line_cache[18][7] ),
    .B2(_09878_),
    .X(_12073_));
 sky130_fd_sc_hd__a221o_1 _16355_ (.A1(\line_cache[17][7] ),
    .A2(_09969_),
    .B1(\line_cache[16][7] ),
    .B2(_09970_),
    .C1(_12073_),
    .X(_12074_));
 sky130_fd_sc_hd__a2111o_1 _16356_ (.A1(\line_cache[20][7] ),
    .A2(_09888_),
    .B1(_12071_),
    .C1(_12072_),
    .D1(_12074_),
    .X(_12075_));
 sky130_fd_sc_hd__a22o_1 _16357_ (.A1(_09796_),
    .A2(\line_cache[33][7] ),
    .B1(\line_cache[34][7] ),
    .B2(_09798_),
    .X(_12076_));
 sky130_fd_sc_hd__a221o_1 _16358_ (.A1(\line_cache[36][7] ),
    .A2(_09777_),
    .B1(\line_cache[35][7] ),
    .B2(_09794_),
    .C1(_12076_),
    .X(_12077_));
 sky130_fd_sc_hd__a22o_1 _16359_ (.A1(_09890_),
    .A2(\line_cache[27][7] ),
    .B1(\line_cache[26][7] ),
    .B2(_09896_),
    .X(_12078_));
 sky130_fd_sc_hd__a221oi_2 _16360_ (.A1(\line_cache[25][7] ),
    .A2(_09892_),
    .B1(\line_cache[24][7] ),
    .B2(_09895_),
    .C1(_12078_),
    .Y(_12079_));
 sky130_fd_sc_hd__a22o_1 _16361_ (.A1(_09903_),
    .A2(\line_cache[29][7] ),
    .B1(\line_cache[28][7] ),
    .B2(_09900_),
    .X(_12080_));
 sky130_fd_sc_hd__a221oi_1 _16362_ (.A1(\line_cache[32][7] ),
    .A2(_09792_),
    .B1(\line_cache[30][7] ),
    .B2(_09905_),
    .C1(_12080_),
    .Y(_12081_));
 sky130_fd_sc_hd__nand2_1 _16363_ (.A(_09773_),
    .B(\line_cache[38][7] ),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_1 _16364_ (.A(_09775_),
    .B(\line_cache[37][7] ),
    .Y(_12083_));
 sky130_fd_sc_hd__nand2_1 _16365_ (.A(_12082_),
    .B(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__a221oi_2 _16366_ (.A1(_09783_),
    .A2(\line_cache[40][7] ),
    .B1(\line_cache[39][7] ),
    .B2(_09780_),
    .C1(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__and4b_1 _16367_ (.A_N(_12077_),
    .B(_12079_),
    .C(_12081_),
    .D(_12085_),
    .X(_12086_));
 sky130_fd_sc_hd__or3b_1 _16368_ (.A(_12070_),
    .B(_12075_),
    .C_N(_12086_),
    .X(_12087_));
 sky130_fd_sc_hd__nor3_2 _16369_ (.A(_12038_),
    .B(_12061_),
    .C(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a22o_1 _16370_ (.A1(_10244_),
    .A2(\line_cache[173][7] ),
    .B1(\line_cache[172][7] ),
    .B2(_10245_),
    .X(_12089_));
 sky130_fd_sc_hd__a221o_1 _16371_ (.A1(\line_cache[175][7] ),
    .A2(_10242_),
    .B1(\line_cache[174][7] ),
    .B2(_10243_),
    .C1(_12089_),
    .X(_12090_));
 sky130_fd_sc_hd__a22o_1 _16372_ (.A1(_10263_),
    .A2(\line_cache[170][7] ),
    .B1(\line_cache[171][7] ),
    .B2(_10262_),
    .X(_12091_));
 sky130_fd_sc_hd__a221o_1 _16373_ (.A1(\line_cache[169][7] ),
    .A2(_10260_),
    .B1(\line_cache[168][7] ),
    .B2(_10261_),
    .C1(_12091_),
    .X(_12092_));
 sky130_fd_sc_hd__a22o_1 _16374_ (.A1(_10256_),
    .A2(\line_cache[160][7] ),
    .B1(\line_cache[161][7] ),
    .B2(_10257_),
    .X(_12093_));
 sky130_fd_sc_hd__and3_1 _16375_ (.A(_10104_),
    .B(_09751_),
    .C(\line_cache[163][7] ),
    .X(_12094_));
 sky130_fd_sc_hd__a22o_1 _16376_ (.A1(_10249_),
    .A2(\line_cache[166][7] ),
    .B1(\line_cache[167][7] ),
    .B2(_10248_),
    .X(_12095_));
 sky130_fd_sc_hd__a221o_1 _16377_ (.A1(\line_cache[165][7] ),
    .A2(_10250_),
    .B1(\line_cache[164][7] ),
    .B2(_10251_),
    .C1(_12095_),
    .X(_12096_));
 sky130_fd_sc_hd__a2111o_1 _16378_ (.A1(\line_cache[162][7] ),
    .A2(_10255_),
    .B1(_12093_),
    .C1(_12094_),
    .D1(_12096_),
    .X(_12097_));
 sky130_fd_sc_hd__nor3_1 _16379_ (.A(_12090_),
    .B(_12092_),
    .C(_12097_),
    .Y(_12098_));
 sky130_fd_sc_hd__a22o_1 _16380_ (.A1(_10272_),
    .A2(\line_cache[189][7] ),
    .B1(\line_cache[188][7] ),
    .B2(_10271_),
    .X(_12099_));
 sky130_fd_sc_hd__a221o_1 _16381_ (.A1(\line_cache[191][7] ),
    .A2(_10269_),
    .B1(\line_cache[190][7] ),
    .B2(_10270_),
    .C1(_12099_),
    .X(_12100_));
 sky130_fd_sc_hd__a22o_1 _16382_ (.A1(_10284_),
    .A2(\line_cache[176][7] ),
    .B1(_10285_),
    .B2(\line_cache[177][7] ),
    .X(_12101_));
 sky130_fd_sc_hd__a221oi_2 _16383_ (.A1(\line_cache[179][7] ),
    .A2(_10282_),
    .B1(\line_cache[178][7] ),
    .B2(_10283_),
    .C1(_12101_),
    .Y(_12102_));
 sky130_fd_sc_hd__and3_1 _16384_ (.A(_10288_),
    .B(_10102_),
    .C(\line_cache[182][7] ),
    .X(_12103_));
 sky130_fd_sc_hd__and3_1 _16385_ (.A(_10288_),
    .B(_10098_),
    .C(\line_cache[181][7] ),
    .X(_12104_));
 sky130_fd_sc_hd__a31o_1 _16386_ (.A1(\line_cache[180][7] ),
    .A2(_10289_),
    .A3(_10106_),
    .B1(_12104_),
    .X(_12105_));
 sky130_fd_sc_hd__a311oi_2 _16387_ (.A1(\line_cache[183][7] ),
    .A2(_10289_),
    .A3(_10061_),
    .B1(_12103_),
    .C1(_12105_),
    .Y(_12106_));
 sky130_fd_sc_hd__a22o_1 _16388_ (.A1(_10277_),
    .A2(\line_cache[184][7] ),
    .B1(\line_cache[185][7] ),
    .B2(_10278_),
    .X(_12107_));
 sky130_fd_sc_hd__a221oi_2 _16389_ (.A1(\line_cache[187][7] ),
    .A2(_10275_),
    .B1(\line_cache[186][7] ),
    .B2(_10276_),
    .C1(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__and4b_1 _16390_ (.A_N(_12100_),
    .B(_12102_),
    .C(_12106_),
    .D(_12108_),
    .X(_12109_));
 sky130_fd_sc_hd__a22o_1 _16391_ (.A1(_10219_),
    .A2(\line_cache[157][7] ),
    .B1(\line_cache[156][7] ),
    .B2(_10220_),
    .X(_12110_));
 sky130_fd_sc_hd__a221o_1 _16392_ (.A1(\line_cache[159][7] ),
    .A2(_10217_),
    .B1(\line_cache[158][7] ),
    .B2(_10218_),
    .C1(_12110_),
    .X(_12111_));
 sky130_fd_sc_hd__a22o_1 _16393_ (.A1(_10238_),
    .A2(\line_cache[154][7] ),
    .B1(\line_cache[155][7] ),
    .B2(_10237_),
    .X(_12112_));
 sky130_fd_sc_hd__a221o_1 _16394_ (.A1(\line_cache[153][7] ),
    .A2(_10235_),
    .B1(\line_cache[152][7] ),
    .B2(_10236_),
    .C1(_12112_),
    .X(_12113_));
 sky130_fd_sc_hd__a22o_1 _16395_ (.A1(_10224_),
    .A2(\line_cache[148][7] ),
    .B1(\line_cache[149][7] ),
    .B2(_10223_),
    .X(_12114_));
 sky130_fd_sc_hd__a22o_1 _16396_ (.A1(_10225_),
    .A2(\line_cache[151][7] ),
    .B1(\line_cache[150][7] ),
    .B2(_10226_),
    .X(_12115_));
 sky130_fd_sc_hd__a22o_1 _16397_ (.A1(_10230_),
    .A2(\line_cache[144][7] ),
    .B1(\line_cache[145][7] ),
    .B2(_10229_),
    .X(_12116_));
 sky130_fd_sc_hd__a22o_1 _16398_ (.A1(_10231_),
    .A2(\line_cache[147][7] ),
    .B1(\line_cache[146][7] ),
    .B2(_10232_),
    .X(_12117_));
 sky130_fd_sc_hd__or4_1 _16399_ (.A(_12114_),
    .B(_12115_),
    .C(_12116_),
    .D(_12117_),
    .X(_12118_));
 sky130_fd_sc_hd__nor3_1 _16400_ (.A(_12111_),
    .B(_12113_),
    .C(_12118_),
    .Y(_12119_));
 sky130_fd_sc_hd__and3_2 _16401_ (.A(_12098_),
    .B(_12109_),
    .C(_12119_),
    .X(_12120_));
 sky130_fd_sc_hd__a22o_1 _16402_ (.A1(_10378_),
    .A2(\line_cache[80][7] ),
    .B1(_10379_),
    .B2(\line_cache[81][7] ),
    .X(_12121_));
 sky130_fd_sc_hd__a221o_1 _16403_ (.A1(\line_cache[83][7] ),
    .A2(_10376_),
    .B1(\line_cache[82][7] ),
    .B2(_10377_),
    .C1(_12121_),
    .X(_12122_));
 sky130_fd_sc_hd__a22o_1 _16404_ (.A1(_10384_),
    .A2(\line_cache[92][7] ),
    .B1(_10385_),
    .B2(\line_cache[93][7] ),
    .X(_12123_));
 sky130_fd_sc_hd__a221o_1 _16405_ (.A1(\line_cache[95][7] ),
    .A2(net136),
    .B1(\line_cache[94][7] ),
    .B2(_10383_),
    .C1(_12123_),
    .X(_12124_));
 sky130_fd_sc_hd__a22o_1 _16406_ (.A1(_10390_),
    .A2(\line_cache[84][7] ),
    .B1(_10391_),
    .B2(\line_cache[85][7] ),
    .X(_12125_));
 sky130_fd_sc_hd__a221o_1 _16407_ (.A1(\line_cache[87][7] ),
    .A2(_10388_),
    .B1(\line_cache[86][7] ),
    .B2(_10389_),
    .C1(_12125_),
    .X(_12126_));
 sky130_fd_sc_hd__a22o_1 _16408_ (.A1(_10396_),
    .A2(\line_cache[88][7] ),
    .B1(_10397_),
    .B2(\line_cache[89][7] ),
    .X(_12127_));
 sky130_fd_sc_hd__a221o_1 _16409_ (.A1(\line_cache[91][7] ),
    .A2(_10394_),
    .B1(\line_cache[90][7] ),
    .B2(_10395_),
    .C1(_12127_),
    .X(_12128_));
 sky130_fd_sc_hd__or4_1 _16410_ (.A(_12122_),
    .B(_12124_),
    .C(_12126_),
    .D(_12128_),
    .X(_12129_));
 sky130_fd_sc_hd__a22o_1 _16411_ (.A1(_10371_),
    .A2(\line_cache[100][7] ),
    .B1(_10372_),
    .B2(\line_cache[101][7] ),
    .X(_12130_));
 sky130_fd_sc_hd__a22o_1 _16412_ (.A1(_10369_),
    .A2(\line_cache[103][7] ),
    .B1(_10370_),
    .B2(\line_cache[102][7] ),
    .X(_12131_));
 sky130_fd_sc_hd__a22o_1 _16413_ (.A1(_10351_),
    .A2(\line_cache[96][7] ),
    .B1(_10352_),
    .B2(\line_cache[97][7] ),
    .X(_12132_));
 sky130_fd_sc_hd__a221o_2 _16414_ (.A1(\line_cache[99][7] ),
    .A2(_10349_),
    .B1(\line_cache[98][7] ),
    .B2(_10348_),
    .C1(_12132_),
    .X(_12133_));
 sky130_fd_sc_hd__and3_1 _16415_ (.A(_10035_),
    .B(\line_cache[107][7] ),
    .C(_10651_),
    .X(_12134_));
 sky130_fd_sc_hd__and3_1 _16416_ (.A(_10176_),
    .B(\line_cache[105][7] ),
    .C(_10651_),
    .X(_12135_));
 sky130_fd_sc_hd__and3_1 _16417_ (.A(_10054_),
    .B(\line_cache[106][7] ),
    .C(_10356_),
    .X(_12136_));
 sky130_fd_sc_hd__and3_1 _16418_ (.A(_10360_),
    .B(\line_cache[104][7] ),
    .C(_10356_),
    .X(_12137_));
 sky130_fd_sc_hd__or4_1 _16419_ (.A(_12134_),
    .B(_12135_),
    .C(_12136_),
    .D(_12137_),
    .X(_12138_));
 sky130_fd_sc_hd__a22o_1 _16420_ (.A1(_10365_),
    .A2(\line_cache[108][7] ),
    .B1(_10366_),
    .B2(\line_cache[109][7] ),
    .X(_12139_));
 sky130_fd_sc_hd__a221o_1 _16421_ (.A1(\line_cache[111][7] ),
    .A2(_10363_),
    .B1(\line_cache[110][7] ),
    .B2(_10364_),
    .C1(_12139_),
    .X(_12140_));
 sky130_fd_sc_hd__or2_1 _16422_ (.A(_12138_),
    .B(_12140_),
    .X(_12141_));
 sky130_fd_sc_hd__or4_1 _16423_ (.A(_12130_),
    .B(_12131_),
    .C(_12133_),
    .D(_12141_),
    .X(_12142_));
 sky130_fd_sc_hd__nor2_1 _16424_ (.A(_12129_),
    .B(_12142_),
    .Y(_12143_));
 sky130_fd_sc_hd__and3_1 _16425_ (.A(_09758_),
    .B(_10031_),
    .C(\line_cache[141][7] ),
    .X(_12144_));
 sky130_fd_sc_hd__a21o_1 _16426_ (.A1(\line_cache[140][7] ),
    .A2(_10336_),
    .B1(_12144_),
    .X(_12145_));
 sky130_fd_sc_hd__a221o_1 _16427_ (.A1(\line_cache[143][7] ),
    .A2(_10334_),
    .B1(\line_cache[142][7] ),
    .B2(_10335_),
    .C1(_12145_),
    .X(_12146_));
 sky130_fd_sc_hd__and3_1 _16428_ (.A(_09758_),
    .B(_10098_),
    .C(\line_cache[133][7] ),
    .X(_12147_));
 sky130_fd_sc_hd__a21o_1 _16429_ (.A1(\line_cache[132][7] ),
    .A2(_10324_),
    .B1(_12147_),
    .X(_12148_));
 sky130_fd_sc_hd__a221o_1 _16430_ (.A1(\line_cache[135][7] ),
    .A2(_10322_),
    .B1(\line_cache[134][7] ),
    .B2(_10323_),
    .C1(_12148_),
    .X(_12149_));
 sky130_fd_sc_hd__and3_1 _16431_ (.A(_10071_),
    .B(\line_cache[128][7] ),
    .C(_09758_),
    .X(_12150_));
 sky130_fd_sc_hd__a21o_1 _16432_ (.A1(\line_cache[129][7] ),
    .A2(_10330_),
    .B1(_12150_),
    .X(_12151_));
 sky130_fd_sc_hd__a221o_1 _16433_ (.A1(\line_cache[131][7] ),
    .A2(_10328_),
    .B1(\line_cache[130][7] ),
    .B2(_10329_),
    .C1(_12151_),
    .X(_12152_));
 sky130_fd_sc_hd__a22o_1 _16434_ (.A1(_10342_),
    .A2(\line_cache[139][7] ),
    .B1(\line_cache[138][7] ),
    .B2(_10343_),
    .X(_12153_));
 sky130_fd_sc_hd__a221o_1 _16435_ (.A1(\line_cache[137][7] ),
    .A2(_10340_),
    .B1(\line_cache[136][7] ),
    .B2(_10341_),
    .C1(_12153_),
    .X(_12154_));
 sky130_fd_sc_hd__or4_1 _16436_ (.A(_12146_),
    .B(_12149_),
    .C(_12152_),
    .D(_12154_),
    .X(_12155_));
 sky130_fd_sc_hd__a22o_1 _16437_ (.A1(_10298_),
    .A2(\line_cache[112][7] ),
    .B1(_10299_),
    .B2(\line_cache[113][7] ),
    .X(_12156_));
 sky130_fd_sc_hd__a221o_1 _16438_ (.A1(\line_cache[115][7] ),
    .A2(_10296_),
    .B1(\line_cache[114][7] ),
    .B2(_10297_),
    .C1(_12156_),
    .X(_12157_));
 sky130_fd_sc_hd__a22o_1 _16439_ (.A1(_10305_),
    .A2(\line_cache[124][7] ),
    .B1(_10306_),
    .B2(\line_cache[125][7] ),
    .X(_12158_));
 sky130_fd_sc_hd__a221o_1 _16440_ (.A1(\line_cache[127][7] ),
    .A2(_10303_),
    .B1(\line_cache[126][7] ),
    .B2(_10304_),
    .C1(_12158_),
    .X(_12159_));
 sky130_fd_sc_hd__a22o_1 _16441_ (.A1(_10311_),
    .A2(\line_cache[116][7] ),
    .B1(_10312_),
    .B2(\line_cache[117][7] ),
    .X(_12160_));
 sky130_fd_sc_hd__a221o_1 _16442_ (.A1(\line_cache[119][7] ),
    .A2(_10309_),
    .B1(\line_cache[118][7] ),
    .B2(_10310_),
    .C1(_12160_),
    .X(_12161_));
 sky130_fd_sc_hd__a22o_1 _16443_ (.A1(_10317_),
    .A2(\line_cache[120][7] ),
    .B1(_10318_),
    .B2(\line_cache[121][7] ),
    .X(_12162_));
 sky130_fd_sc_hd__a221o_1 _16444_ (.A1(\line_cache[123][7] ),
    .A2(_10315_),
    .B1(\line_cache[122][7] ),
    .B2(_10316_),
    .C1(_12162_),
    .X(_12163_));
 sky130_fd_sc_hd__or4_1 _16445_ (.A(_12157_),
    .B(_12159_),
    .C(_12161_),
    .D(_12163_),
    .X(_12164_));
 sky130_fd_sc_hd__nor2_1 _16446_ (.A(_12155_),
    .B(_12164_),
    .Y(_12165_));
 sky130_fd_sc_hd__and3_1 _16447_ (.A(_12120_),
    .B(_12143_),
    .C(_12165_),
    .X(_12166_));
 sky130_fd_sc_hd__nand3_1 _16448_ (.A(_12025_),
    .B(_12088_),
    .C(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__o21ba_2 _16449_ (.A1(_11918_),
    .A2(_12167_),
    .B1_N(_08979_),
    .X(_12168_));
 sky130_fd_sc_hd__buf_6 _16450_ (.A(_12168_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_16 _16451_ (.A(net66),
    .X(_12169_));
 sky130_fd_sc_hd__clkbuf_16 _16452_ (.A(_12169_),
    .X(_12170_));
 sky130_fd_sc_hd__nand2_8 _16453_ (.A(net3921),
    .B(net3982),
    .Y(_12171_));
 sky130_fd_sc_hd__nand2_1 _16454_ (.A(net3995),
    .B(net3381),
    .Y(_12172_));
 sky130_fd_sc_hd__inv_2 _16455_ (.A(_12172_),
    .Y(_12173_));
 sky130_fd_sc_hd__nor2_2 _16456_ (.A(\line_cache_idx[7] ),
    .B(\line_cache_idx[6] ),
    .Y(_12174_));
 sky130_fd_sc_hd__nand2_2 _16457_ (.A(_12173_),
    .B(_12174_),
    .Y(_12175_));
 sky130_fd_sc_hd__nor2_1 _16458_ (.A(_12171_),
    .B(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__buf_6 _16459_ (.A(_09070_),
    .X(_12177_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(_12176_),
    .B(_12177_),
    .Y(_12178_));
 sky130_fd_sc_hd__buf_4 _16461_ (.A(_12178_),
    .X(_12179_));
 sky130_fd_sc_hd__buf_8 _16462_ (.A(_09125_),
    .X(_12180_));
 sky130_fd_sc_hd__clkbuf_8 _16463_ (.A(_12180_),
    .X(_12181_));
 sky130_fd_sc_hd__buf_4 _16464_ (.A(_12178_),
    .X(_12182_));
 sky130_fd_sc_hd__clkbuf_8 _16465_ (.A(net50),
    .X(_12183_));
 sky130_fd_sc_hd__inv_8 _16466_ (.A(_12183_),
    .Y(_12184_));
 sky130_fd_sc_hd__buf_8 _16467_ (.A(_12184_),
    .X(_12185_));
 sky130_fd_sc_hd__nand2_1 _16468_ (.A(_12182_),
    .B(_12185_),
    .Y(_12186_));
 sky130_fd_sc_hd__o211a_1 _16469_ (.A1(_12170_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12186_),
    .X(_12187_));
 sky130_fd_sc_hd__nand2_4 _16470_ (.A(net75),
    .B(_09106_),
    .Y(_12188_));
 sky130_fd_sc_hd__nand2_8 _16471_ (.A(_12188_),
    .B(net49),
    .Y(_12189_));
 sky130_fd_sc_hd__buf_12 _16472_ (.A(_12189_),
    .X(_12190_));
 sky130_fd_sc_hd__a21bo_1 _16473_ (.A1(_12178_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_12191_));
 sky130_fd_sc_hd__clkbuf_8 _16474_ (.A(_12191_),
    .X(_12192_));
 sky130_fd_sc_hd__mux2_1 _16475_ (.A0(_12187_),
    .A1(net3757),
    .S(_12192_),
    .X(_12193_));
 sky130_fd_sc_hd__clkbuf_1 _16476_ (.A(_12193_),
    .X(_00012_));
 sky130_fd_sc_hd__buf_12 _16477_ (.A(net67),
    .X(_12194_));
 sky130_fd_sc_hd__clkbuf_16 _16478_ (.A(_12194_),
    .X(_12195_));
 sky130_fd_sc_hd__clkbuf_8 _16479_ (.A(net61),
    .X(_12196_));
 sky130_fd_sc_hd__inv_12 _16480_ (.A(_12196_),
    .Y(_12197_));
 sky130_fd_sc_hd__clkbuf_16 _16481_ (.A(_12197_),
    .X(_12198_));
 sky130_fd_sc_hd__nand2_1 _16482_ (.A(_12182_),
    .B(_12198_),
    .Y(_12199_));
 sky130_fd_sc_hd__o211a_1 _16483_ (.A1(_12195_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12199_),
    .X(_12200_));
 sky130_fd_sc_hd__mux2_1 _16484_ (.A0(_12200_),
    .A1(net3810),
    .S(_12192_),
    .X(_12201_));
 sky130_fd_sc_hd__clkbuf_1 _16485_ (.A(_12201_),
    .X(_00013_));
 sky130_fd_sc_hd__clkbuf_16 _16486_ (.A(net68),
    .X(_12202_));
 sky130_fd_sc_hd__buf_12 _16487_ (.A(_12202_),
    .X(_12203_));
 sky130_fd_sc_hd__buf_6 _16488_ (.A(net72),
    .X(_12204_));
 sky130_fd_sc_hd__inv_12 _16489_ (.A(_12204_),
    .Y(_12205_));
 sky130_fd_sc_hd__clkbuf_16 _16490_ (.A(_12205_),
    .X(_12206_));
 sky130_fd_sc_hd__nand2_1 _16491_ (.A(_12182_),
    .B(_12206_),
    .Y(_12207_));
 sky130_fd_sc_hd__o211a_1 _16492_ (.A1(_12203_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12207_),
    .X(_12208_));
 sky130_fd_sc_hd__mux2_1 _16493_ (.A0(_12208_),
    .A1(net3643),
    .S(_12192_),
    .X(_12209_));
 sky130_fd_sc_hd__clkbuf_1 _16494_ (.A(_12209_),
    .X(_00014_));
 sky130_fd_sc_hd__clkbuf_16 _16495_ (.A(net69),
    .X(_12210_));
 sky130_fd_sc_hd__clkbuf_16 _16496_ (.A(_12210_),
    .X(_12211_));
 sky130_fd_sc_hd__buf_8 _16497_ (.A(net76),
    .X(_12212_));
 sky130_fd_sc_hd__inv_12 _16498_ (.A(_12212_),
    .Y(_12213_));
 sky130_fd_sc_hd__clkbuf_16 _16499_ (.A(_12213_),
    .X(_12214_));
 sky130_fd_sc_hd__nand2_1 _16500_ (.A(_12182_),
    .B(_12214_),
    .Y(_12215_));
 sky130_fd_sc_hd__o211a_1 _16501_ (.A1(_12211_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12215_),
    .X(_12216_));
 sky130_fd_sc_hd__mux2_1 _16502_ (.A0(_12216_),
    .A1(net3685),
    .S(_12192_),
    .X(_12217_));
 sky130_fd_sc_hd__clkbuf_1 _16503_ (.A(_12217_),
    .X(_00015_));
 sky130_fd_sc_hd__clkbuf_16 _16504_ (.A(net70),
    .X(_12218_));
 sky130_fd_sc_hd__buf_12 _16505_ (.A(_12218_),
    .X(_12219_));
 sky130_fd_sc_hd__buf_6 _16506_ (.A(net77),
    .X(_12220_));
 sky130_fd_sc_hd__inv_12 _16507_ (.A(_12220_),
    .Y(_12221_));
 sky130_fd_sc_hd__buf_12 _16508_ (.A(_12221_),
    .X(_12222_));
 sky130_fd_sc_hd__nand2_1 _16509_ (.A(_12182_),
    .B(_12222_),
    .Y(_12223_));
 sky130_fd_sc_hd__o211a_1 _16510_ (.A1(_12219_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12223_),
    .X(_12224_));
 sky130_fd_sc_hd__mux2_1 _16511_ (.A0(_12224_),
    .A1(net3623),
    .S(_12192_),
    .X(_12225_));
 sky130_fd_sc_hd__clkbuf_1 _16512_ (.A(_12225_),
    .X(_00016_));
 sky130_fd_sc_hd__clkbuf_16 _16513_ (.A(net71),
    .X(_12226_));
 sky130_fd_sc_hd__clkbuf_16 _16514_ (.A(_12226_),
    .X(_12227_));
 sky130_fd_sc_hd__buf_6 _16515_ (.A(net78),
    .X(_12228_));
 sky130_fd_sc_hd__inv_8 _16516_ (.A(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__clkbuf_16 _16517_ (.A(_12229_),
    .X(_12230_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(_12182_),
    .B(_12230_),
    .Y(_12231_));
 sky130_fd_sc_hd__o211a_1 _16519_ (.A1(_12227_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12231_),
    .X(_12232_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(_12232_),
    .A1(net3762),
    .S(_12192_),
    .X(_12233_));
 sky130_fd_sc_hd__clkbuf_1 _16521_ (.A(_12233_),
    .X(_00017_));
 sky130_fd_sc_hd__clkbuf_16 _16522_ (.A(net73),
    .X(_12234_));
 sky130_fd_sc_hd__clkbuf_16 _16523_ (.A(_12234_),
    .X(_12235_));
 sky130_fd_sc_hd__clkbuf_8 _16524_ (.A(net79),
    .X(_12236_));
 sky130_fd_sc_hd__inv_8 _16525_ (.A(_12236_),
    .Y(_12237_));
 sky130_fd_sc_hd__buf_12 _16526_ (.A(_12237_),
    .X(_12238_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(_12182_),
    .B(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__o211a_1 _16528_ (.A1(_12235_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12239_),
    .X(_12240_));
 sky130_fd_sc_hd__mux2_1 _16529_ (.A0(_12240_),
    .A1(net3771),
    .S(_12192_),
    .X(_12241_));
 sky130_fd_sc_hd__clkbuf_1 _16530_ (.A(_12241_),
    .X(_00018_));
 sky130_fd_sc_hd__clkbuf_16 _16531_ (.A(net74),
    .X(_12242_));
 sky130_fd_sc_hd__clkbuf_16 _16532_ (.A(_12242_),
    .X(_12243_));
 sky130_fd_sc_hd__clkbuf_8 _16533_ (.A(net80),
    .X(_12244_));
 sky130_fd_sc_hd__inv_8 _16534_ (.A(_12244_),
    .Y(_12245_));
 sky130_fd_sc_hd__clkbuf_16 _16535_ (.A(_12245_),
    .X(_12246_));
 sky130_fd_sc_hd__nand2_1 _16536_ (.A(_12182_),
    .B(_12246_),
    .Y(_12247_));
 sky130_fd_sc_hd__o211a_1 _16537_ (.A1(_12243_),
    .A2(_12179_),
    .B1(_12181_),
    .C1(_12247_),
    .X(_12248_));
 sky130_fd_sc_hd__mux2_1 _16538_ (.A0(_12248_),
    .A1(net3692),
    .S(_12192_),
    .X(_12249_));
 sky130_fd_sc_hd__clkbuf_1 _16539_ (.A(_12249_),
    .X(_00019_));
 sky130_fd_sc_hd__nor2_1 _16540_ (.A(net88),
    .B(net89),
    .Y(_12250_));
 sky130_fd_sc_hd__inv_2 _16541_ (.A(net91),
    .Y(_12251_));
 sky130_fd_sc_hd__and3_1 _16542_ (.A(_12250_),
    .B(net90),
    .C(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__buf_4 _16543_ (.A(_12252_),
    .X(_12253_));
 sky130_fd_sc_hd__or3b_2 _16544_ (.A(net90),
    .B(_12251_),
    .C_N(_12250_),
    .X(_12254_));
 sky130_fd_sc_hd__clkinv_4 _16545_ (.A(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__nor2_4 _16546_ (.A(_12253_),
    .B(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__a22o_1 _16547_ (.A1(net32),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net33),
    .X(_12257_));
 sky130_fd_sc_hd__a21o_1 _16548_ (.A1(net31),
    .A2(_12256_),
    .B1(_12257_),
    .X(_12258_));
 sky130_fd_sc_hd__inv_2 _16549_ (.A(net88),
    .Y(_12259_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(net90),
    .B(net91),
    .Y(_12260_));
 sky130_fd_sc_hd__inv_2 _16551_ (.A(_12256_),
    .Y(_12261_));
 sky130_fd_sc_hd__a31o_1 _16552_ (.A1(_12259_),
    .A2(net89),
    .A3(_12260_),
    .B1(_12261_),
    .X(_12262_));
 sky130_fd_sc_hd__nand2_1 _16553_ (.A(_12262_),
    .B(_09057_),
    .Y(_12263_));
 sky130_fd_sc_hd__clkbuf_8 _16554_ (.A(_12263_),
    .X(_12264_));
 sky130_fd_sc_hd__mux2_1 _16555_ (.A0(_12258_),
    .A1(net3880),
    .S(_12264_),
    .X(_12265_));
 sky130_fd_sc_hd__clkbuf_1 _16556_ (.A(_12265_),
    .X(_00020_));
 sky130_fd_sc_hd__a22o_1 _16557_ (.A1(net33),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net34),
    .X(_12266_));
 sky130_fd_sc_hd__a21o_1 _16558_ (.A1(net32),
    .A2(_12256_),
    .B1(_12266_),
    .X(_12267_));
 sky130_fd_sc_hd__mux2_1 _16559_ (.A0(_12267_),
    .A1(net3853),
    .S(_12264_),
    .X(_12268_));
 sky130_fd_sc_hd__clkbuf_1 _16560_ (.A(_12268_),
    .X(_00021_));
 sky130_fd_sc_hd__inv_2 _16561_ (.A(net33),
    .Y(_12269_));
 sky130_fd_sc_hd__nor2_1 _16562_ (.A(_12269_),
    .B(_12261_),
    .Y(_12270_));
 sky130_fd_sc_hd__a221o_1 _16563_ (.A1(net34),
    .A2(_12253_),
    .B1(net35),
    .B2(_12255_),
    .C1(_12270_),
    .X(_12271_));
 sky130_fd_sc_hd__mux2_1 _16564_ (.A0(_12271_),
    .A1(net3758),
    .S(_12264_),
    .X(_12272_));
 sky130_fd_sc_hd__clkbuf_1 _16565_ (.A(_12272_),
    .X(_00022_));
 sky130_fd_sc_hd__a22o_1 _16566_ (.A1(net35),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net36),
    .X(_12273_));
 sky130_fd_sc_hd__a21o_1 _16567_ (.A1(net34),
    .A2(_12256_),
    .B1(_12273_),
    .X(_12274_));
 sky130_fd_sc_hd__mux2_1 _16568_ (.A0(_12274_),
    .A1(net3780),
    .S(_12264_),
    .X(_12275_));
 sky130_fd_sc_hd__clkbuf_1 _16569_ (.A(_12275_),
    .X(_00023_));
 sky130_fd_sc_hd__inv_2 _16570_ (.A(net35),
    .Y(_12276_));
 sky130_fd_sc_hd__nor2_1 _16571_ (.A(_12276_),
    .B(_12261_),
    .Y(_12277_));
 sky130_fd_sc_hd__a221o_1 _16572_ (.A1(net36),
    .A2(_12253_),
    .B1(net37),
    .B2(_12255_),
    .C1(_12277_),
    .X(_12278_));
 sky130_fd_sc_hd__mux2_1 _16573_ (.A0(_12278_),
    .A1(net3747),
    .S(_12264_),
    .X(_12279_));
 sky130_fd_sc_hd__clkbuf_1 _16574_ (.A(_12279_),
    .X(_00024_));
 sky130_fd_sc_hd__a22o_1 _16575_ (.A1(net37),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net38),
    .X(_12280_));
 sky130_fd_sc_hd__a21o_1 _16576_ (.A1(net36),
    .A2(_12256_),
    .B1(_12280_),
    .X(_12281_));
 sky130_fd_sc_hd__mux2_1 _16577_ (.A0(_12281_),
    .A1(net3704),
    .S(_12264_),
    .X(_12282_));
 sky130_fd_sc_hd__clkbuf_1 _16578_ (.A(_12282_),
    .X(_00025_));
 sky130_fd_sc_hd__a22o_1 _16579_ (.A1(net38),
    .A2(_12253_),
    .B1(_12256_),
    .B2(net37),
    .X(_12283_));
 sky130_fd_sc_hd__mux2_1 _16580_ (.A0(_12283_),
    .A1(net3820),
    .S(_12264_),
    .X(_12284_));
 sky130_fd_sc_hd__clkbuf_1 _16581_ (.A(_12284_),
    .X(_00026_));
 sky130_fd_sc_hd__inv_2 _16582_ (.A(net38),
    .Y(_12285_));
 sky130_fd_sc_hd__nor2_1 _16583_ (.A(_12285_),
    .B(_12261_),
    .Y(_12286_));
 sky130_fd_sc_hd__mux2_1 _16584_ (.A0(_12286_),
    .A1(net3863),
    .S(_12264_),
    .X(_12287_));
 sky130_fd_sc_hd__clkbuf_1 _16585_ (.A(_12287_),
    .X(_00027_));
 sky130_fd_sc_hd__inv_2 _16586_ (.A(net3982),
    .Y(_12288_));
 sky130_fd_sc_hd__inv_6 _16587_ (.A(_09109_),
    .Y(_12289_));
 sky130_fd_sc_hd__buf_12 _16588_ (.A(_12289_),
    .X(_12290_));
 sky130_fd_sc_hd__or3_1 _16589_ (.A(net3982),
    .B(_12290_),
    .C(_09105_),
    .X(_12291_));
 sky130_fd_sc_hd__o21ai_1 _16590_ (.A1(_12288_),
    .A2(_09110_),
    .B1(net3983),
    .Y(_00028_));
 sky130_fd_sc_hd__nand2_8 _16591_ (.A(_12288_),
    .B(net3921),
    .Y(_12292_));
 sky130_fd_sc_hd__nand2_8 _16592_ (.A(_09081_),
    .B(\line_cache_idx[2] ),
    .Y(_12293_));
 sky130_fd_sc_hd__a21oi_1 _16593_ (.A1(_12292_),
    .A2(_12293_),
    .B1(_12290_),
    .Y(_12294_));
 sky130_fd_sc_hd__a22o_1 _16594_ (.A1(net3921),
    .A2(_12290_),
    .B1(_09112_),
    .B2(_12294_),
    .X(_00029_));
 sky130_fd_sc_hd__or3_1 _16595_ (.A(_09090_),
    .B(_12171_),
    .C(_12290_),
    .X(_12295_));
 sky130_fd_sc_hd__inv_2 _16596_ (.A(_12171_),
    .Y(_12296_));
 sky130_fd_sc_hd__a21o_1 _16597_ (.A1(_09110_),
    .A2(_12296_),
    .B1(net3995),
    .X(_12297_));
 sky130_fd_sc_hd__and3_1 _16598_ (.A(_09111_),
    .B(_12295_),
    .C(_12297_),
    .X(_12298_));
 sky130_fd_sc_hd__clkbuf_1 _16599_ (.A(_12298_),
    .X(_00030_));
 sky130_fd_sc_hd__o21ai_1 _16600_ (.A1(_09090_),
    .A2(_12171_),
    .B1(_09092_),
    .Y(_12299_));
 sky130_fd_sc_hd__nor2_1 _16601_ (.A(_12171_),
    .B(_12172_),
    .Y(_12300_));
 sky130_fd_sc_hd__inv_2 _16602_ (.A(_12300_),
    .Y(_12301_));
 sky130_fd_sc_hd__and3_1 _16603_ (.A(_12299_),
    .B(_12301_),
    .C(_09110_),
    .X(_12302_));
 sky130_fd_sc_hd__a22o_1 _16604_ (.A1(net3381),
    .A2(_12290_),
    .B1(_09112_),
    .B2(_12302_),
    .X(_00031_));
 sky130_fd_sc_hd__inv_2 _16605_ (.A(net4001),
    .Y(_12303_));
 sky130_fd_sc_hd__or3_1 _16606_ (.A(_12303_),
    .B(_12290_),
    .C(_12301_),
    .X(_12304_));
 sky130_fd_sc_hd__a21o_1 _16607_ (.A1(_12300_),
    .A2(_09110_),
    .B1(net4001),
    .X(_12305_));
 sky130_fd_sc_hd__and3_1 _16608_ (.A(_09111_),
    .B(_12304_),
    .C(_12305_),
    .X(_12306_));
 sky130_fd_sc_hd__clkbuf_1 _16609_ (.A(_12306_),
    .X(_00032_));
 sky130_fd_sc_hd__a21o_1 _16610_ (.A1(_12300_),
    .A2(\line_cache_idx[6] ),
    .B1(net3913),
    .X(_12307_));
 sky130_fd_sc_hd__nand2_2 _16611_ (.A(net3913),
    .B(\line_cache_idx[6] ),
    .Y(_12308_));
 sky130_fd_sc_hd__nor2_2 _16612_ (.A(_12308_),
    .B(_12301_),
    .Y(_12309_));
 sky130_fd_sc_hd__nor2_1 _16613_ (.A(_12290_),
    .B(_12309_),
    .Y(_12310_));
 sky130_fd_sc_hd__a32o_1 _16614_ (.A1(_09112_),
    .A2(_12307_),
    .A3(_12310_),
    .B1(net3913),
    .B2(_12290_),
    .X(_00033_));
 sky130_fd_sc_hd__nor2_2 _16615_ (.A(_12172_),
    .B(_12308_),
    .Y(_12311_));
 sky130_fd_sc_hd__a31o_1 _16616_ (.A1(_12311_),
    .A2(_09110_),
    .A3(_12296_),
    .B1(_12177_),
    .X(_12312_));
 sky130_fd_sc_hd__clkbuf_16 _16617_ (.A(_09071_),
    .X(_12313_));
 sky130_fd_sc_hd__or3b_1 _16618_ (.A(_12313_),
    .B(_12289_),
    .C_N(_12309_),
    .X(_12314_));
 sky130_fd_sc_hd__and3_1 _16619_ (.A(_09111_),
    .B(_12312_),
    .C(_12314_),
    .X(_12315_));
 sky130_fd_sc_hd__clkbuf_1 _16620_ (.A(_12315_),
    .X(_00034_));
 sky130_fd_sc_hd__or2_1 _16621_ (.A(_09077_),
    .B(_12314_),
    .X(_12316_));
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(_12314_),
    .B(_09077_),
    .Y(_12317_));
 sky130_fd_sc_hd__and3_1 _16623_ (.A(_09111_),
    .B(_12316_),
    .C(_12317_),
    .X(_12318_));
 sky130_fd_sc_hd__clkbuf_1 _16624_ (.A(_12318_),
    .X(_00035_));
 sky130_fd_sc_hd__nor2_1 _16625_ (.A(net2003),
    .B(net3829),
    .Y(_12319_));
 sky130_fd_sc_hd__inv_2 _16626_ (.A(net3749),
    .Y(_12320_));
 sky130_fd_sc_hd__inv_2 _16627_ (.A(net3804),
    .Y(_12321_));
 sky130_fd_sc_hd__and3_1 _16628_ (.A(_12319_),
    .B(_12320_),
    .C(_12321_),
    .X(_12322_));
 sky130_fd_sc_hd__nor2_1 _16629_ (.A(net2057),
    .B(net2028),
    .Y(_12323_));
 sky130_fd_sc_hd__nand2_1 _16630_ (.A(_12322_),
    .B(_12323_),
    .Y(_12324_));
 sky130_fd_sc_hd__or4_2 _16631_ (.A(net3777),
    .B(net2497),
    .C(net3836),
    .D(net3451),
    .X(_12325_));
 sky130_fd_sc_hd__o21ai_4 _16632_ (.A1(_12324_),
    .A2(_12325_),
    .B1(\fb_read_state[2] ),
    .Y(_12326_));
 sky130_fd_sc_hd__nand2_1 _16633_ (.A(_09107_),
    .B(\fb_read_state[2] ),
    .Y(_12327_));
 sky130_fd_sc_hd__a21oi_4 _16634_ (.A1(_12327_),
    .A2(_12188_),
    .B1(_09056_),
    .Y(_12328_));
 sky130_fd_sc_hd__nand2_2 _16635_ (.A(_12326_),
    .B(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__inv_2 _16636_ (.A(_12329_),
    .Y(_12330_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(_12330_),
    .B(_09106_),
    .Y(_12331_));
 sky130_fd_sc_hd__inv_2 _16638_ (.A(_12331_),
    .Y(_12332_));
 sky130_fd_sc_hd__buf_4 _16639_ (.A(_12330_),
    .X(_12333_));
 sky130_fd_sc_hd__nand2_1 _16640_ (.A(_12333_),
    .B(net2561),
    .Y(_12334_));
 sky130_fd_sc_hd__o21a_1 _16641_ (.A1(net2561),
    .A2(_12332_),
    .B1(_12334_),
    .X(_00036_));
 sky130_fd_sc_hd__nand2_1 _16642_ (.A(net2561),
    .B(net3900),
    .Y(_12335_));
 sky130_fd_sc_hd__or2_1 _16643_ (.A(net2561),
    .B(net3900),
    .X(_12336_));
 sky130_fd_sc_hd__buf_4 _16644_ (.A(_12329_),
    .X(_12337_));
 sky130_fd_sc_hd__and2_1 _16645_ (.A(_12337_),
    .B(net3900),
    .X(_12338_));
 sky130_fd_sc_hd__a41o_1 _16646_ (.A1(_12333_),
    .A2(_09106_),
    .A3(_12335_),
    .A4(_12336_),
    .B1(_12338_),
    .X(_00037_));
 sky130_fd_sc_hd__or2_1 _16647_ (.A(_12335_),
    .B(_12337_),
    .X(_12339_));
 sky130_fd_sc_hd__inv_2 _16648_ (.A(net3557),
    .Y(_12340_));
 sky130_fd_sc_hd__nand2_4 _16649_ (.A(_12330_),
    .B(_09107_),
    .Y(_12341_));
 sky130_fd_sc_hd__inv_2 _16650_ (.A(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__or2_1 _16651_ (.A(_12340_),
    .B(_12335_),
    .X(_12343_));
 sky130_fd_sc_hd__or2_1 _16652_ (.A(_12343_),
    .B(_12329_),
    .X(_12344_));
 sky130_fd_sc_hd__inv_2 _16653_ (.A(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__a211oi_1 _16654_ (.A1(_12339_),
    .A2(_12340_),
    .B1(_12342_),
    .C1(_12345_),
    .Y(_00038_));
 sky130_fd_sc_hd__nor2b_1 _16655_ (.A(_12343_),
    .B_N(net3764),
    .Y(_12346_));
 sky130_fd_sc_hd__nand2_1 _16656_ (.A(_12333_),
    .B(_12346_),
    .Y(_12347_));
 sky130_fd_sc_hd__o211a_1 _16657_ (.A1(net3764),
    .A2(_12345_),
    .B1(_12341_),
    .C1(_12347_),
    .X(_00039_));
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(_12346_),
    .B(net3854),
    .Y(_12348_));
 sky130_fd_sc_hd__a31o_1 _16659_ (.A1(_12326_),
    .A2(_12328_),
    .A3(_12346_),
    .B1(net3854),
    .X(_12349_));
 sky130_fd_sc_hd__o211a_1 _16660_ (.A1(_12337_),
    .A2(_12348_),
    .B1(_12341_),
    .C1(net3855),
    .X(_00040_));
 sky130_fd_sc_hd__a31o_1 _16661_ (.A1(_12333_),
    .A2(net3854),
    .A3(_12346_),
    .B1(net3987),
    .X(_12350_));
 sky130_fd_sc_hd__nand2b_1 _16662_ (.A_N(_12348_),
    .B(net3987),
    .Y(_12351_));
 sky130_fd_sc_hd__or2_1 _16663_ (.A(_12351_),
    .B(_12337_),
    .X(_12352_));
 sky130_fd_sc_hd__and3_1 _16664_ (.A(_12350_),
    .B(_12341_),
    .C(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__clkbuf_1 _16665_ (.A(_12353_),
    .X(_00041_));
 sky130_fd_sc_hd__inv_2 _16666_ (.A(net3624),
    .Y(_12354_));
 sky130_fd_sc_hd__or2_1 _16667_ (.A(_12354_),
    .B(_12351_),
    .X(_12355_));
 sky130_fd_sc_hd__inv_2 _16668_ (.A(_12355_),
    .Y(_12356_));
 sky130_fd_sc_hd__nand2_1 _16669_ (.A(_12330_),
    .B(_12356_),
    .Y(_12357_));
 sky130_fd_sc_hd__inv_2 _16670_ (.A(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__a211oi_1 _16671_ (.A1(_12352_),
    .A2(_12354_),
    .B1(_12342_),
    .C1(_12358_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_1 _16672_ (.A(_12356_),
    .B(net2750),
    .Y(_12359_));
 sky130_fd_sc_hd__inv_2 _16673_ (.A(_12359_),
    .Y(_12360_));
 sky130_fd_sc_hd__nand2_1 _16674_ (.A(_12360_),
    .B(_12330_),
    .Y(_12361_));
 sky130_fd_sc_hd__o211a_1 _16675_ (.A1(net2750),
    .A2(_12358_),
    .B1(_12341_),
    .C1(_12361_),
    .X(_00043_));
 sky130_fd_sc_hd__inv_2 _16676_ (.A(net3618),
    .Y(_12362_));
 sky130_fd_sc_hd__nor2_1 _16677_ (.A(_12362_),
    .B(_12361_),
    .Y(_12363_));
 sky130_fd_sc_hd__or2_1 _16678_ (.A(_12342_),
    .B(_12363_),
    .X(_12364_));
 sky130_fd_sc_hd__a21oi_1 _16679_ (.A1(_12362_),
    .A2(_12361_),
    .B1(_12364_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand2_1 _16680_ (.A(net3618),
    .B(net3768),
    .Y(_12365_));
 sky130_fd_sc_hd__nor2_1 _16681_ (.A(_12365_),
    .B(_12359_),
    .Y(_12366_));
 sky130_fd_sc_hd__nand2_1 _16682_ (.A(_12366_),
    .B(_12330_),
    .Y(_12367_));
 sky130_fd_sc_hd__o211a_1 _16683_ (.A1(net3768),
    .A2(_12363_),
    .B1(_12341_),
    .C1(_12367_),
    .X(_00045_));
 sky130_fd_sc_hd__inv_2 _16684_ (.A(net3821),
    .Y(_12368_));
 sky130_fd_sc_hd__nor2_1 _16685_ (.A(_12368_),
    .B(_12367_),
    .Y(_12369_));
 sky130_fd_sc_hd__or2_1 _16686_ (.A(_12342_),
    .B(_12369_),
    .X(_12370_));
 sky130_fd_sc_hd__a21oi_1 _16687_ (.A1(_12368_),
    .A2(_12367_),
    .B1(_12370_),
    .Y(_00046_));
 sky130_fd_sc_hd__inv_2 _16688_ (.A(net3497),
    .Y(_12371_));
 sky130_fd_sc_hd__inv_2 _16689_ (.A(_12366_),
    .Y(_12372_));
 sky130_fd_sc_hd__or4_1 _16690_ (.A(_12368_),
    .B(_12371_),
    .C(_12329_),
    .D(_12372_),
    .X(_12373_));
 sky130_fd_sc_hd__o211a_1 _16691_ (.A1(net3497),
    .A2(_12369_),
    .B1(_12341_),
    .C1(_12373_),
    .X(_00047_));
 sky130_fd_sc_hd__inv_2 _16692_ (.A(net3790),
    .Y(_12374_));
 sky130_fd_sc_hd__or4_1 _16693_ (.A(_12368_),
    .B(_12371_),
    .C(_12374_),
    .D(_12372_),
    .X(_12375_));
 sky130_fd_sc_hd__nor2_1 _16694_ (.A(_12337_),
    .B(_12375_),
    .Y(_12376_));
 sky130_fd_sc_hd__a211oi_1 _16695_ (.A1(_12373_),
    .A2(_12374_),
    .B1(_12342_),
    .C1(_12376_),
    .Y(_00048_));
 sky130_fd_sc_hd__nor2b_1 _16696_ (.A(_12375_),
    .B_N(net3494),
    .Y(_12377_));
 sky130_fd_sc_hd__nand2_1 _16697_ (.A(_12377_),
    .B(_12330_),
    .Y(_12378_));
 sky130_fd_sc_hd__o211a_1 _16698_ (.A1(net3494),
    .A2(_12376_),
    .B1(_12341_),
    .C1(_12378_),
    .X(_00049_));
 sky130_fd_sc_hd__inv_2 _16699_ (.A(net3792),
    .Y(_12379_));
 sky130_fd_sc_hd__nor2_1 _16700_ (.A(_12379_),
    .B(_12378_),
    .Y(_12380_));
 sky130_fd_sc_hd__or2_1 _16701_ (.A(_12342_),
    .B(_12380_),
    .X(_12381_));
 sky130_fd_sc_hd__a21oi_1 _16702_ (.A1(_12379_),
    .A2(_12378_),
    .B1(_12381_),
    .Y(_00050_));
 sky130_fd_sc_hd__inv_2 _16703_ (.A(net3660),
    .Y(_12382_));
 sky130_fd_sc_hd__or3b_1 _16704_ (.A(_12379_),
    .B(_12382_),
    .C_N(_12377_),
    .X(_12383_));
 sky130_fd_sc_hd__o221a_1 _16705_ (.A1(net3660),
    .A2(_12380_),
    .B1(_12337_),
    .B2(_12383_),
    .C1(_12341_),
    .X(_00051_));
 sky130_fd_sc_hd__or3_1 _16706_ (.A(net3846),
    .B(_12337_),
    .C(_12383_),
    .X(_12384_));
 sky130_fd_sc_hd__o21ai_1 _16707_ (.A1(_12337_),
    .A2(_12383_),
    .B1(net3846),
    .Y(_12385_));
 sky130_fd_sc_hd__a21oi_1 _16708_ (.A1(net3847),
    .A2(_12385_),
    .B1(_12342_),
    .Y(_00052_));
 sky130_fd_sc_hd__nand2_1 _16709_ (.A(net3790),
    .B(net106),
    .Y(_12386_));
 sky130_fd_sc_hd__or3_1 _16710_ (.A(_12368_),
    .B(_12371_),
    .C(_12365_),
    .X(_12387_));
 sky130_fd_sc_hd__or4_1 _16711_ (.A(_12379_),
    .B(_12382_),
    .C(_12386_),
    .D(_12387_),
    .X(_12388_));
 sky130_fd_sc_hd__nor2_1 _16712_ (.A(_12359_),
    .B(_12388_),
    .Y(_12389_));
 sky130_fd_sc_hd__a21o_1 _16713_ (.A1(_12389_),
    .A2(net109),
    .B1(net2009),
    .X(_12390_));
 sky130_fd_sc_hd__nand2_1 _16714_ (.A(net3846),
    .B(net2009),
    .Y(_12391_));
 sky130_fd_sc_hd__inv_2 _16715_ (.A(_12391_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand2_1 _16716_ (.A(_12389_),
    .B(_12392_),
    .Y(_12393_));
 sky130_fd_sc_hd__a32o_1 _16717_ (.A1(_12390_),
    .A2(_12332_),
    .A3(_12393_),
    .B1(net2009),
    .B2(_12337_),
    .X(_00053_));
 sky130_fd_sc_hd__inv_2 _16718_ (.A(net3996),
    .Y(_12394_));
 sky130_fd_sc_hd__or3_1 _16719_ (.A(_12394_),
    .B(_12337_),
    .C(_12393_),
    .X(_12395_));
 sky130_fd_sc_hd__o21ai_1 _16720_ (.A1(_12337_),
    .A2(_12393_),
    .B1(_12394_),
    .Y(_12396_));
 sky130_fd_sc_hd__and3_1 _16721_ (.A(_12395_),
    .B(_12341_),
    .C(_12396_),
    .X(_12397_));
 sky130_fd_sc_hd__clkbuf_1 _16722_ (.A(_12397_),
    .X(_00054_));
 sky130_fd_sc_hd__inv_2 _16723_ (.A(net3016),
    .Y(_12398_));
 sky130_fd_sc_hd__or2_1 _16724_ (.A(_12394_),
    .B(_12393_),
    .X(_12399_));
 sky130_fd_sc_hd__nor2_1 _16725_ (.A(_12398_),
    .B(_12399_),
    .Y(_12400_));
 sky130_fd_sc_hd__nor2_1 _16726_ (.A(_12331_),
    .B(_12400_),
    .Y(_12401_));
 sky130_fd_sc_hd__nand2_1 _16727_ (.A(_12399_),
    .B(_12398_),
    .Y(_12402_));
 sky130_fd_sc_hd__a22o_1 _16728_ (.A1(net3016),
    .A2(_12337_),
    .B1(_12401_),
    .B2(_12402_),
    .X(_00055_));
 sky130_fd_sc_hd__a21oi_1 _16729_ (.A1(_12400_),
    .A2(_12333_),
    .B1(net3841),
    .Y(_12403_));
 sky130_fd_sc_hd__a31o_1 _16730_ (.A1(_12400_),
    .A2(net3841),
    .A3(_12333_),
    .B1(_12342_),
    .X(_12404_));
 sky130_fd_sc_hd__nor2_1 _16731_ (.A(net3842),
    .B(_12404_),
    .Y(_00056_));
 sky130_fd_sc_hd__and3_1 _16732_ (.A(_12400_),
    .B(net3841),
    .C(net2021),
    .X(_12405_));
 sky130_fd_sc_hd__and3_1 _16733_ (.A(_12392_),
    .B(net111),
    .C(net3016),
    .X(_12406_));
 sky130_fd_sc_hd__a31o_1 _16734_ (.A1(_12389_),
    .A2(net113),
    .A3(_12406_),
    .B1(net2021),
    .X(_12407_));
 sky130_fd_sc_hd__or3b_1 _16735_ (.A(_12331_),
    .B(_12405_),
    .C_N(_12407_),
    .X(_12408_));
 sky130_fd_sc_hd__a21bo_1 _16736_ (.A1(net2021),
    .A2(_12337_),
    .B1_N(_12408_),
    .X(_00057_));
 sky130_fd_sc_hd__a21oi_1 _16737_ (.A1(_12405_),
    .A2(_12333_),
    .B1(net3860),
    .Y(_12409_));
 sky130_fd_sc_hd__and3_1 _16738_ (.A(_12405_),
    .B(net3860),
    .C(_12333_),
    .X(_12410_));
 sky130_fd_sc_hd__nor3_1 _16739_ (.A(_12342_),
    .B(net3861),
    .C(_12410_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand3_1 _16740_ (.A(_12405_),
    .B(net115),
    .C(net3607),
    .Y(_12411_));
 sky130_fd_sc_hd__o221a_1 _16741_ (.A1(_12337_),
    .A2(_12411_),
    .B1(net3607),
    .B2(_12410_),
    .C1(_12341_),
    .X(_00059_));
 sky130_fd_sc_hd__inv_2 _16742_ (.A(net3950),
    .Y(_12412_));
 sky130_fd_sc_hd__and4_1 _16743_ (.A(net3841),
    .B(net2021),
    .C(net3860),
    .D(net3607),
    .X(_12413_));
 sky130_fd_sc_hd__and2_1 _16744_ (.A(_12413_),
    .B(_12406_),
    .X(_12414_));
 sky130_fd_sc_hd__nand2_1 _16745_ (.A(_12389_),
    .B(_12414_),
    .Y(_12415_));
 sky130_fd_sc_hd__or2_1 _16746_ (.A(_12412_),
    .B(_12415_),
    .X(_12416_));
 sky130_fd_sc_hd__nand2_1 _16747_ (.A(_12415_),
    .B(_12412_),
    .Y(_12417_));
 sky130_fd_sc_hd__nor2_1 _16748_ (.A(_12412_),
    .B(_12333_),
    .Y(_12418_));
 sky130_fd_sc_hd__a41o_1 _16749_ (.A1(_12416_),
    .A2(_12417_),
    .A3(_09106_),
    .A4(_12333_),
    .B1(_12418_),
    .X(_00060_));
 sky130_fd_sc_hd__inv_2 _16750_ (.A(net2017),
    .Y(_12419_));
 sky130_fd_sc_hd__or3_1 _16751_ (.A(_12412_),
    .B(_12419_),
    .C(_12411_),
    .X(_12420_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(_12416_),
    .B(_12419_),
    .Y(_12421_));
 sky130_fd_sc_hd__a32o_1 _16753_ (.A1(_12420_),
    .A2(_12332_),
    .A3(_12421_),
    .B1(net2017),
    .B2(_12337_),
    .X(_00061_));
 sky130_fd_sc_hd__inv_2 _16754_ (.A(net3975),
    .Y(_12422_));
 sky130_fd_sc_hd__nand2_1 _16755_ (.A(net3950),
    .B(net2017),
    .Y(_12423_));
 sky130_fd_sc_hd__or2_1 _16756_ (.A(_12423_),
    .B(_12415_),
    .X(_12424_));
 sky130_fd_sc_hd__or2_1 _16757_ (.A(_12422_),
    .B(_12424_),
    .X(_12425_));
 sky130_fd_sc_hd__nand2_1 _16758_ (.A(_12424_),
    .B(_12422_),
    .Y(_12426_));
 sky130_fd_sc_hd__nor2_1 _16759_ (.A(_12422_),
    .B(_12333_),
    .Y(_12427_));
 sky130_fd_sc_hd__a41o_1 _16760_ (.A1(_12425_),
    .A2(_12426_),
    .A3(_09106_),
    .A4(_12333_),
    .B1(_12427_),
    .X(_00062_));
 sky130_fd_sc_hd__inv_2 _16761_ (.A(net2007),
    .Y(_12428_));
 sky130_fd_sc_hd__or3_1 _16762_ (.A(_12422_),
    .B(_12428_),
    .C(_12420_),
    .X(_12429_));
 sky130_fd_sc_hd__nand2_1 _16763_ (.A(_12425_),
    .B(_12428_),
    .Y(_12430_));
 sky130_fd_sc_hd__a32o_1 _16764_ (.A1(_12429_),
    .A2(_12332_),
    .A3(_12430_),
    .B1(net2007),
    .B2(_12337_),
    .X(_00063_));
 sky130_fd_sc_hd__inv_2 _16765_ (.A(net3956),
    .Y(_12431_));
 sky130_fd_sc_hd__or4_1 _16766_ (.A(_12422_),
    .B(_12428_),
    .C(_12423_),
    .D(_12415_),
    .X(_12432_));
 sky130_fd_sc_hd__or2_1 _16767_ (.A(_12431_),
    .B(_12432_),
    .X(_12433_));
 sky130_fd_sc_hd__nand2_1 _16768_ (.A(_12432_),
    .B(_12431_),
    .Y(_12434_));
 sky130_fd_sc_hd__nor2_1 _16769_ (.A(_12431_),
    .B(_12333_),
    .Y(_12435_));
 sky130_fd_sc_hd__a41o_1 _16770_ (.A1(_12433_),
    .A2(_12434_),
    .A3(_09106_),
    .A4(_12333_),
    .B1(_12435_),
    .X(_00064_));
 sky130_fd_sc_hd__inv_2 _16771_ (.A(net3962),
    .Y(_12436_));
 sky130_fd_sc_hd__or2_1 _16772_ (.A(_12436_),
    .B(_12433_),
    .X(_12437_));
 sky130_fd_sc_hd__nand2_1 _16773_ (.A(_12433_),
    .B(_12436_),
    .Y(_12438_));
 sky130_fd_sc_hd__nor2_1 _16774_ (.A(_12436_),
    .B(_12333_),
    .Y(_12439_));
 sky130_fd_sc_hd__a41o_1 _16775_ (.A1(_12437_),
    .A2(_09106_),
    .A3(_12438_),
    .A4(_12333_),
    .B1(_12439_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _16776_ (.A0(net84),
    .A1(net3952),
    .S(_09516_),
    .X(_12440_));
 sky130_fd_sc_hd__clkbuf_1 _16777_ (.A(_12440_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _16778_ (.A0(net85),
    .A1(net3866),
    .S(_09516_),
    .X(_12441_));
 sky130_fd_sc_hd__clkbuf_1 _16779_ (.A(_12441_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _16780_ (.A0(net86),
    .A1(net3756),
    .S(_09516_),
    .X(_12442_));
 sky130_fd_sc_hd__clkbuf_1 _16781_ (.A(_12442_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _16782_ (.A0(net87),
    .A1(net3891),
    .S(_09516_),
    .X(_12443_));
 sky130_fd_sc_hd__clkbuf_1 _16783_ (.A(_12443_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _16784_ (.A0(net88),
    .A1(net3907),
    .S(_09516_),
    .X(_12444_));
 sky130_fd_sc_hd__clkbuf_1 _16785_ (.A(_12444_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _16786_ (.A0(net89),
    .A1(net3735),
    .S(_09516_),
    .X(_12445_));
 sky130_fd_sc_hd__clkbuf_1 _16787_ (.A(_12445_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _16788_ (.A0(net90),
    .A1(net3763),
    .S(_09516_),
    .X(_12446_));
 sky130_fd_sc_hd__clkbuf_1 _16789_ (.A(_12446_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _16790_ (.A0(net91),
    .A1(net3738),
    .S(_09516_),
    .X(_12447_));
 sky130_fd_sc_hd__clkbuf_1 _16791_ (.A(_12447_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _16792_ (.A0(net1),
    .A1(net3923),
    .S(_09516_),
    .X(_12448_));
 sky130_fd_sc_hd__clkbuf_1 _16793_ (.A(_12448_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _16794_ (.A0(net2),
    .A1(net3942),
    .S(_09516_),
    .X(_12449_));
 sky130_fd_sc_hd__clkbuf_1 _16795_ (.A(_12449_),
    .X(_00075_));
 sky130_fd_sc_hd__clkbuf_8 _16796_ (.A(_09126_),
    .X(_12450_));
 sky130_fd_sc_hd__mux2_1 _16797_ (.A0(net3),
    .A1(net3895),
    .S(_12450_),
    .X(_12451_));
 sky130_fd_sc_hd__clkbuf_1 _16798_ (.A(_12451_),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _16799_ (.A0(net4),
    .A1(net3961),
    .S(_12450_),
    .X(_12452_));
 sky130_fd_sc_hd__clkbuf_1 _16800_ (.A(_12452_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _16801_ (.A0(net5),
    .A1(net3896),
    .S(_12450_),
    .X(_12453_));
 sky130_fd_sc_hd__clkbuf_1 _16802_ (.A(_12453_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _16803_ (.A0(net6),
    .A1(net3940),
    .S(_12450_),
    .X(_12454_));
 sky130_fd_sc_hd__clkbuf_1 _16804_ (.A(_12454_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _16805_ (.A0(net7),
    .A1(net3928),
    .S(_12450_),
    .X(_12455_));
 sky130_fd_sc_hd__clkbuf_1 _16806_ (.A(_12455_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _16807_ (.A0(net8),
    .A1(net3844),
    .S(_12450_),
    .X(_12456_));
 sky130_fd_sc_hd__clkbuf_1 _16808_ (.A(_12456_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _16809_ (.A0(net9),
    .A1(net3911),
    .S(_12450_),
    .X(_12457_));
 sky130_fd_sc_hd__clkbuf_1 _16810_ (.A(_12457_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _16811_ (.A0(net10),
    .A1(net3870),
    .S(_12450_),
    .X(_12458_));
 sky130_fd_sc_hd__clkbuf_1 _16812_ (.A(_12458_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _16813_ (.A0(net18),
    .A1(net3698),
    .S(_12450_),
    .X(_12459_));
 sky130_fd_sc_hd__clkbuf_1 _16814_ (.A(_12459_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _16815_ (.A0(net19),
    .A1(net3877),
    .S(_12450_),
    .X(_12460_));
 sky130_fd_sc_hd__clkbuf_1 _16816_ (.A(_12460_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _16817_ (.A0(net20),
    .A1(net3832),
    .S(_12450_),
    .X(_12461_));
 sky130_fd_sc_hd__clkbuf_1 _16818_ (.A(_12461_),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _16819_ (.A0(net21),
    .A1(net3887),
    .S(_12450_),
    .X(_12462_));
 sky130_fd_sc_hd__clkbuf_1 _16820_ (.A(_12462_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _16821_ (.A0(net22),
    .A1(net3707),
    .S(_12450_),
    .X(_12463_));
 sky130_fd_sc_hd__clkbuf_1 _16822_ (.A(_12463_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _16823_ (.A0(net23),
    .A1(net3701),
    .S(_12450_),
    .X(_12464_));
 sky130_fd_sc_hd__clkbuf_1 _16824_ (.A(_12464_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _16825_ (.A0(net24),
    .A1(net3934),
    .S(_12450_),
    .X(_12465_));
 sky130_fd_sc_hd__clkbuf_1 _16826_ (.A(_12465_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _16827_ (.A0(net25),
    .A1(net3926),
    .S(_12450_),
    .X(_12466_));
 sky130_fd_sc_hd__clkbuf_1 _16828_ (.A(_12466_),
    .X(_00091_));
 sky130_fd_sc_hd__buf_6 _16829_ (.A(_09126_),
    .X(_12467_));
 sky130_fd_sc_hd__mux2_1 _16830_ (.A0(net26),
    .A1(net3893),
    .S(_12467_),
    .X(_12468_));
 sky130_fd_sc_hd__clkbuf_1 _16831_ (.A(_12468_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _16832_ (.A0(net27),
    .A1(net3834),
    .S(_12467_),
    .X(_12469_));
 sky130_fd_sc_hd__clkbuf_1 _16833_ (.A(_12469_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _16834_ (.A0(net28),
    .A1(net3857),
    .S(_12467_),
    .X(_12470_));
 sky130_fd_sc_hd__clkbuf_1 _16835_ (.A(_12470_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _16836_ (.A0(net29),
    .A1(net3918),
    .S(_12467_),
    .X(_12471_));
 sky130_fd_sc_hd__clkbuf_1 _16837_ (.A(_12471_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _16838_ (.A0(net11),
    .A1(net3816),
    .S(_12467_),
    .X(_12472_));
 sky130_fd_sc_hd__clkbuf_1 _16839_ (.A(_12472_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _16840_ (.A0(net12),
    .A1(net3932),
    .S(_12467_),
    .X(_12473_));
 sky130_fd_sc_hd__clkbuf_1 _16841_ (.A(_12473_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _16842_ (.A0(net13),
    .A1(net3953),
    .S(_12467_),
    .X(_12474_));
 sky130_fd_sc_hd__clkbuf_1 _16843_ (.A(_12474_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _16844_ (.A0(net14),
    .A1(net3881),
    .S(_12467_),
    .X(_12475_));
 sky130_fd_sc_hd__clkbuf_1 _16845_ (.A(_12475_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _16846_ (.A0(net15),
    .A1(net3894),
    .S(_12467_),
    .X(_12476_));
 sky130_fd_sc_hd__clkbuf_1 _16847_ (.A(_12476_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _16848_ (.A0(net16),
    .A1(net3884),
    .S(_12467_),
    .X(_12477_));
 sky130_fd_sc_hd__clkbuf_1 _16849_ (.A(_12477_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _16850_ (.A0(net17),
    .A1(net3935),
    .S(_12467_),
    .X(_12478_));
 sky130_fd_sc_hd__clkbuf_1 _16851_ (.A(_12478_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _16852_ (.A0(net30),
    .A1(net3927),
    .S(_12467_),
    .X(_12479_));
 sky130_fd_sc_hd__clkbuf_1 _16853_ (.A(_12479_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _16854_ (.A0(net31),
    .A1(net3835),
    .S(_12467_),
    .X(_12480_));
 sky130_fd_sc_hd__clkbuf_1 _16855_ (.A(_12480_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _16856_ (.A0(net32),
    .A1(net3850),
    .S(_12467_),
    .X(_12481_));
 sky130_fd_sc_hd__clkbuf_1 _16857_ (.A(_12481_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _16858_ (.A0(net33),
    .A1(net3949),
    .S(_12467_),
    .X(_12482_));
 sky130_fd_sc_hd__clkbuf_1 _16859_ (.A(_12482_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _16860_ (.A0(net34),
    .A1(net3938),
    .S(_12467_),
    .X(_12483_));
 sky130_fd_sc_hd__clkbuf_1 _16861_ (.A(_12483_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _16862_ (.A0(net35),
    .A1(net3908),
    .S(_09127_),
    .X(_12484_));
 sky130_fd_sc_hd__clkbuf_1 _16863_ (.A(_12484_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _16864_ (.A0(net36),
    .A1(net3954),
    .S(_09127_),
    .X(_12485_));
 sky130_fd_sc_hd__clkbuf_1 _16865_ (.A(_12485_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _16866_ (.A0(net37),
    .A1(net3906),
    .S(_09127_),
    .X(_12486_));
 sky130_fd_sc_hd__clkbuf_1 _16867_ (.A(_12486_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _16868_ (.A0(net38),
    .A1(net3815),
    .S(_09127_),
    .X(_12487_));
 sky130_fd_sc_hd__clkbuf_1 _16869_ (.A(_12487_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _16870_ (.A0(net43),
    .A1(net3595),
    .S(_09127_),
    .X(_12488_));
 sky130_fd_sc_hd__clkbuf_1 _16871_ (.A(_12488_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _16872_ (.A0(net44),
    .A1(net3852),
    .S(_09127_),
    .X(_12489_));
 sky130_fd_sc_hd__clkbuf_1 _16873_ (.A(_12489_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _16874_ (.A0(net45),
    .A1(net3838),
    .S(_09127_),
    .X(_12490_));
 sky130_fd_sc_hd__clkbuf_1 _16875_ (.A(_12490_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _16876_ (.A0(net46),
    .A1(net3486),
    .S(_09127_),
    .X(_12491_));
 sky130_fd_sc_hd__clkbuf_1 _16877_ (.A(_12491_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _16878_ (.A0(net47),
    .A1(net3876),
    .S(_09127_),
    .X(_12492_));
 sky130_fd_sc_hd__clkbuf_1 _16879_ (.A(_12492_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _16880_ (.A0(net48),
    .A1(net3905),
    .S(_09127_),
    .X(_12493_));
 sky130_fd_sc_hd__clkbuf_1 _16881_ (.A(_12493_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _16882_ (.A0(net39),
    .A1(net3939),
    .S(_09127_),
    .X(_12494_));
 sky130_fd_sc_hd__clkbuf_1 _16883_ (.A(_12494_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _16884_ (.A0(net40),
    .A1(net3904),
    .S(_09127_),
    .X(_12495_));
 sky130_fd_sc_hd__clkbuf_1 _16885_ (.A(_12495_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _16886_ (.A0(net41),
    .A1(net3964),
    .S(_09127_),
    .X(_12496_));
 sky130_fd_sc_hd__clkbuf_1 _16887_ (.A(_12496_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _16888_ (.A0(net42),
    .A1(net3897),
    .S(_09127_),
    .X(_12497_));
 sky130_fd_sc_hd__clkbuf_1 _16889_ (.A(_12497_),
    .X(_00121_));
 sky130_fd_sc_hd__a22o_1 _16890_ (.A1(net3),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net4),
    .X(_12498_));
 sky130_fd_sc_hd__a21o_1 _16891_ (.A1(net2),
    .A2(_12256_),
    .B1(_12498_),
    .X(_12499_));
 sky130_fd_sc_hd__mux2_1 _16892_ (.A0(_12499_),
    .A1(net3929),
    .S(_12264_),
    .X(_12500_));
 sky130_fd_sc_hd__clkbuf_1 _16893_ (.A(_12500_),
    .X(_00122_));
 sky130_fd_sc_hd__a22o_1 _16894_ (.A1(net4),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net5),
    .X(_12501_));
 sky130_fd_sc_hd__a21o_1 _16895_ (.A1(net3),
    .A2(_12256_),
    .B1(_12501_),
    .X(_12502_));
 sky130_fd_sc_hd__mux2_1 _16896_ (.A0(_12502_),
    .A1(net3910),
    .S(_12264_),
    .X(_12503_));
 sky130_fd_sc_hd__clkbuf_1 _16897_ (.A(_12503_),
    .X(_00123_));
 sky130_fd_sc_hd__a22o_1 _16898_ (.A1(net5),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net6),
    .X(_12504_));
 sky130_fd_sc_hd__a21o_1 _16899_ (.A1(net4),
    .A2(_12256_),
    .B1(_12504_),
    .X(_12505_));
 sky130_fd_sc_hd__mux2_1 _16900_ (.A0(_12505_),
    .A1(net3974),
    .S(_12264_),
    .X(_12506_));
 sky130_fd_sc_hd__clkbuf_1 _16901_ (.A(_12506_),
    .X(_00124_));
 sky130_fd_sc_hd__a22o_1 _16902_ (.A1(net6),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net7),
    .X(_12507_));
 sky130_fd_sc_hd__a21o_1 _16903_ (.A1(net5),
    .A2(_12256_),
    .B1(_12507_),
    .X(_12508_));
 sky130_fd_sc_hd__mux2_1 _16904_ (.A0(_12508_),
    .A1(net3931),
    .S(_12264_),
    .X(_12509_));
 sky130_fd_sc_hd__clkbuf_1 _16905_ (.A(_12509_),
    .X(_00125_));
 sky130_fd_sc_hd__a22o_1 _16906_ (.A1(net7),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net8),
    .X(_12510_));
 sky130_fd_sc_hd__a21o_1 _16907_ (.A1(net6),
    .A2(_12256_),
    .B1(_12510_),
    .X(_12511_));
 sky130_fd_sc_hd__mux2_1 _16908_ (.A0(_12511_),
    .A1(net3945),
    .S(_12264_),
    .X(_12512_));
 sky130_fd_sc_hd__clkbuf_1 _16909_ (.A(_12512_),
    .X(_00126_));
 sky130_fd_sc_hd__a22o_1 _16910_ (.A1(net8),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net9),
    .X(_12513_));
 sky130_fd_sc_hd__a21o_1 _16911_ (.A1(net7),
    .A2(_12256_),
    .B1(_12513_),
    .X(_12514_));
 sky130_fd_sc_hd__mux2_1 _16912_ (.A0(_12514_),
    .A1(net3967),
    .S(_12264_),
    .X(_12515_));
 sky130_fd_sc_hd__clkbuf_1 _16913_ (.A(_12515_),
    .X(_00127_));
 sky130_fd_sc_hd__a22o_1 _16914_ (.A1(net9),
    .A2(_12253_),
    .B1(_12255_),
    .B2(net10),
    .X(_12516_));
 sky130_fd_sc_hd__a21o_1 _16915_ (.A1(net8),
    .A2(_12256_),
    .B1(_12516_),
    .X(_12517_));
 sky130_fd_sc_hd__mux2_1 _16916_ (.A0(_12517_),
    .A1(net3970),
    .S(_12264_),
    .X(_12518_));
 sky130_fd_sc_hd__clkbuf_1 _16917_ (.A(_12518_),
    .X(_00128_));
 sky130_fd_sc_hd__a22o_1 _16918_ (.A1(net10),
    .A2(_12253_),
    .B1(_12256_),
    .B2(net9),
    .X(_12519_));
 sky130_fd_sc_hd__mux2_1 _16919_ (.A0(_12519_),
    .A1(net3966),
    .S(_12264_),
    .X(_12520_));
 sky130_fd_sc_hd__clkbuf_1 _16920_ (.A(_12520_),
    .X(_00129_));
 sky130_fd_sc_hd__and2_1 _16921_ (.A(_12256_),
    .B(net10),
    .X(_12521_));
 sky130_fd_sc_hd__mux2_1 _16922_ (.A0(_12521_),
    .A1(net3971),
    .S(_12263_),
    .X(_12522_));
 sky130_fd_sc_hd__clkbuf_1 _16923_ (.A(_12522_),
    .X(_00130_));
 sky130_fd_sc_hd__inv_2 _16924_ (.A(\base_h_bporch[6] ),
    .Y(_12523_));
 sky130_fd_sc_hd__nand2_1 _16925_ (.A(_09297_),
    .B(_12523_),
    .Y(_12524_));
 sky130_fd_sc_hd__nand3_2 _16926_ (.A(_09257_),
    .B(\base_h_bporch[6] ),
    .C(_09296_),
    .Y(_12525_));
 sky130_fd_sc_hd__nand2_1 _16927_ (.A(_12524_),
    .B(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__nor2_1 _16928_ (.A(_09259_),
    .B(_12526_),
    .Y(_12527_));
 sky130_fd_sc_hd__inv_2 _16929_ (.A(\base_h_bporch[1] ),
    .Y(_12528_));
 sky130_fd_sc_hd__nand2_1 _16930_ (.A(_09282_),
    .B(_12528_),
    .Y(_12529_));
 sky130_fd_sc_hd__nand3_1 _16931_ (.A(_09211_),
    .B(_09281_),
    .C(\base_h_bporch[1] ),
    .Y(_12530_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(_09286_),
    .B(\base_h_bporch[0] ),
    .Y(_12531_));
 sky130_fd_sc_hd__inv_2 _16933_ (.A(_12531_),
    .Y(_12532_));
 sky130_fd_sc_hd__nand3_1 _16934_ (.A(_12529_),
    .B(_12530_),
    .C(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__nand2_1 _16935_ (.A(_12533_),
    .B(_12530_),
    .Y(_12534_));
 sky130_fd_sc_hd__nand3_1 _16936_ (.A(_09221_),
    .B(_09273_),
    .C(\base_h_bporch[2] ),
    .Y(_12535_));
 sky130_fd_sc_hd__inv_2 _16937_ (.A(\base_h_bporch[2] ),
    .Y(_12536_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(_09274_),
    .B(_12536_),
    .Y(_12537_));
 sky130_fd_sc_hd__nand3_1 _16939_ (.A(_12534_),
    .B(_12535_),
    .C(_12537_),
    .Y(_12538_));
 sky130_fd_sc_hd__nand2_1 _16940_ (.A(_12538_),
    .B(_12535_),
    .Y(_12539_));
 sky130_fd_sc_hd__inv_2 _16941_ (.A(\base_h_bporch[3] ),
    .Y(_12540_));
 sky130_fd_sc_hd__nand2_1 _16942_ (.A(_09278_),
    .B(_12540_),
    .Y(_12541_));
 sky130_fd_sc_hd__nand2_1 _16943_ (.A(_12539_),
    .B(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__or2_1 _16944_ (.A(_12540_),
    .B(_09278_),
    .X(_12543_));
 sky130_fd_sc_hd__nand2_1 _16945_ (.A(_12542_),
    .B(_12543_),
    .Y(_12544_));
 sky130_fd_sc_hd__inv_2 _16946_ (.A(\base_h_bporch[5] ),
    .Y(_12545_));
 sky130_fd_sc_hd__nand2_1 _16947_ (.A(_09267_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__nand3_2 _16948_ (.A(_09264_),
    .B(_09266_),
    .C(\base_h_bporch[5] ),
    .Y(_12547_));
 sky130_fd_sc_hd__inv_2 _16949_ (.A(\base_h_bporch[4] ),
    .Y(_12548_));
 sky130_fd_sc_hd__nand2_1 _16950_ (.A(_09269_),
    .B(_12548_),
    .Y(_12549_));
 sky130_fd_sc_hd__nand3_2 _16951_ (.A(_09262_),
    .B(_09268_),
    .C(\base_h_bporch[4] ),
    .Y(_12550_));
 sky130_fd_sc_hd__nand2_1 _16952_ (.A(_12549_),
    .B(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__inv_2 _16953_ (.A(_12551_),
    .Y(_12552_));
 sky130_fd_sc_hd__nand3_1 _16954_ (.A(_12546_),
    .B(_12547_),
    .C(_12552_),
    .Y(_12553_));
 sky130_fd_sc_hd__inv_2 _16955_ (.A(_12553_),
    .Y(_12554_));
 sky130_fd_sc_hd__nand3_1 _16956_ (.A(_12527_),
    .B(_12544_),
    .C(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__nor2_1 _16957_ (.A(_12525_),
    .B(_09259_),
    .Y(_12556_));
 sky130_fd_sc_hd__inv_2 _16958_ (.A(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__inv_2 _16959_ (.A(_12550_),
    .Y(_12558_));
 sky130_fd_sc_hd__nand3_1 _16960_ (.A(_12546_),
    .B(_12547_),
    .C(_12558_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand2_1 _16961_ (.A(_12559_),
    .B(_12547_),
    .Y(_12560_));
 sky130_fd_sc_hd__nand2_1 _16962_ (.A(_12527_),
    .B(_12560_),
    .Y(_12561_));
 sky130_fd_sc_hd__nand3_1 _16963_ (.A(_12555_),
    .B(_12557_),
    .C(_12561_),
    .Y(_12562_));
 sky130_fd_sc_hd__nand2_1 _16964_ (.A(_12562_),
    .B(_09247_),
    .Y(_12563_));
 sky130_fd_sc_hd__nand2_1 _16965_ (.A(_12563_),
    .B(_09250_),
    .Y(_12564_));
 sky130_fd_sc_hd__nand3_1 _16966_ (.A(_12562_),
    .B(_09251_),
    .C(_09247_),
    .Y(_12565_));
 sky130_fd_sc_hd__nand2_1 _16967_ (.A(_12564_),
    .B(_12565_),
    .Y(_12566_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(_12552_),
    .B(_12544_),
    .Y(_12567_));
 sky130_fd_sc_hd__nand2_1 _16969_ (.A(_12567_),
    .B(_12550_),
    .Y(_12568_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(_09267_),
    .B(\base_h_bporch[5] ),
    .Y(_12569_));
 sky130_fd_sc_hd__nand3_1 _16971_ (.A(_09264_),
    .B(_09266_),
    .C(_12545_),
    .Y(_12570_));
 sky130_fd_sc_hd__nand2_1 _16972_ (.A(_12569_),
    .B(_12570_),
    .Y(_12571_));
 sky130_fd_sc_hd__nand2_1 _16973_ (.A(_12568_),
    .B(_12571_),
    .Y(_12572_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(_12572_),
    .B(_12547_),
    .Y(_12573_));
 sky130_fd_sc_hd__inv_2 _16975_ (.A(_12526_),
    .Y(_12574_));
 sky130_fd_sc_hd__nand2_1 _16976_ (.A(_12573_),
    .B(_12574_),
    .Y(_12575_));
 sky130_fd_sc_hd__nand3_1 _16977_ (.A(_12572_),
    .B(_12547_),
    .C(_12526_),
    .Y(_12576_));
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(_12575_),
    .B(_12576_),
    .Y(_12577_));
 sky130_fd_sc_hd__nand2_1 _16979_ (.A(_12546_),
    .B(_12547_),
    .Y(_12578_));
 sky130_fd_sc_hd__nand3_1 _16980_ (.A(_12578_),
    .B(_12550_),
    .C(_12567_),
    .Y(_12579_));
 sky130_fd_sc_hd__nand2_1 _16981_ (.A(_12579_),
    .B(_12572_),
    .Y(_12580_));
 sky130_fd_sc_hd__nand3_1 _16982_ (.A(_12551_),
    .B(_12543_),
    .C(_12542_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand2_1 _16983_ (.A(_12581_),
    .B(_12567_),
    .Y(_12582_));
 sky130_fd_sc_hd__a21boi_1 _16984_ (.A1(_12534_),
    .A2(_12537_),
    .B1_N(_12535_),
    .Y(_12583_));
 sky130_fd_sc_hd__nand3_1 _16985_ (.A(_09275_),
    .B(_09277_),
    .C(_12540_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand2_1 _16986_ (.A(_09278_),
    .B(\base_h_bporch[3] ),
    .Y(_12585_));
 sky130_fd_sc_hd__nand3_1 _16987_ (.A(_12583_),
    .B(_12584_),
    .C(_12585_),
    .Y(_12586_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(_12585_),
    .B(_12584_),
    .Y(_12587_));
 sky130_fd_sc_hd__nand2_1 _16989_ (.A(_12587_),
    .B(_12539_),
    .Y(_12588_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(_12586_),
    .B(_12588_),
    .Y(_12589_));
 sky130_fd_sc_hd__inv_2 _16991_ (.A(_12534_),
    .Y(_12590_));
 sky130_fd_sc_hd__nand2_1 _16992_ (.A(_12537_),
    .B(_12535_),
    .Y(_12591_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(_12590_),
    .B(_12591_),
    .Y(_12592_));
 sky130_fd_sc_hd__nand2_1 _16994_ (.A(_12538_),
    .B(_12592_),
    .Y(_12593_));
 sky130_fd_sc_hd__nand2_1 _16995_ (.A(_12529_),
    .B(_12530_),
    .Y(_12594_));
 sky130_fd_sc_hd__nand2_1 _16996_ (.A(_12594_),
    .B(_12531_),
    .Y(_12595_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(_12595_),
    .B(_12533_),
    .Y(_12596_));
 sky130_fd_sc_hd__or2_1 _16998_ (.A(\base_h_bporch[0] ),
    .B(_09286_),
    .X(_12597_));
 sky130_fd_sc_hd__nand2_1 _16999_ (.A(_12597_),
    .B(_12531_),
    .Y(_12598_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_12596_),
    .B(_12598_),
    .Y(_12599_));
 sky130_fd_sc_hd__inv_2 _17001_ (.A(_12599_),
    .Y(_12600_));
 sky130_fd_sc_hd__nand2_1 _17002_ (.A(_12593_),
    .B(_12600_),
    .Y(_12601_));
 sky130_fd_sc_hd__inv_2 _17003_ (.A(_12601_),
    .Y(_12602_));
 sky130_fd_sc_hd__nand2_2 _17004_ (.A(_12589_),
    .B(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__inv_2 _17005_ (.A(_12603_),
    .Y(_12604_));
 sky130_fd_sc_hd__nand2_1 _17006_ (.A(_12582_),
    .B(_12604_),
    .Y(_12605_));
 sky130_fd_sc_hd__inv_2 _17007_ (.A(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__nand2_1 _17008_ (.A(_12580_),
    .B(_12606_),
    .Y(_12607_));
 sky130_fd_sc_hd__inv_2 _17009_ (.A(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(_12577_),
    .B(_12608_),
    .Y(_12609_));
 sky130_fd_sc_hd__nand2_1 _17011_ (.A(_12575_),
    .B(_12525_),
    .Y(_12610_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(_12610_),
    .B(_09259_),
    .Y(_12611_));
 sky130_fd_sc_hd__nand3_1 _17013_ (.A(_12575_),
    .B(_09260_),
    .C(_12525_),
    .Y(_12612_));
 sky130_fd_sc_hd__nand2_1 _17014_ (.A(_12611_),
    .B(_12612_),
    .Y(_12613_));
 sky130_fd_sc_hd__nor2_1 _17015_ (.A(_12609_),
    .B(_12613_),
    .Y(_12614_));
 sky130_fd_sc_hd__a21oi_1 _17016_ (.A1(_12527_),
    .A2(_12560_),
    .B1(_12556_),
    .Y(_12615_));
 sky130_fd_sc_hd__nand3_1 _17017_ (.A(_12615_),
    .B(_09246_),
    .C(_12555_),
    .Y(_12616_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(_12563_),
    .B(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__nand3_1 _17019_ (.A(_12566_),
    .B(_12614_),
    .C(_12617_),
    .Y(_12618_));
 sky130_fd_sc_hd__inv_2 _17020_ (.A(_12609_),
    .Y(_12619_));
 sky130_fd_sc_hd__nand2_1 _17021_ (.A(_12613_),
    .B(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__nand2_1 _17022_ (.A(_12610_),
    .B(_09260_),
    .Y(_12621_));
 sky130_fd_sc_hd__nand3_1 _17023_ (.A(_12575_),
    .B(_09259_),
    .C(_12525_),
    .Y(_12622_));
 sky130_fd_sc_hd__nand2_1 _17024_ (.A(_12621_),
    .B(_12622_),
    .Y(_12623_));
 sky130_fd_sc_hd__nand2_1 _17025_ (.A(_12623_),
    .B(_12609_),
    .Y(_12624_));
 sky130_fd_sc_hd__nand2_1 _17026_ (.A(_12620_),
    .B(_12624_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand2_1 _17027_ (.A(_12625_),
    .B(net3968),
    .Y(_12626_));
 sky130_fd_sc_hd__nand2_1 _17028_ (.A(_12618_),
    .B(_12626_),
    .Y(_12627_));
 sky130_fd_sc_hd__nand3_1 _17029_ (.A(_12620_),
    .B(_12624_),
    .C(_08874_),
    .Y(_12628_));
 sky130_fd_sc_hd__nand3_1 _17030_ (.A(_12603_),
    .B(_12581_),
    .C(_12567_),
    .Y(_12629_));
 sky130_fd_sc_hd__a21oi_1 _17031_ (.A1(_12605_),
    .A2(_12629_),
    .B1(\base_h_counter[4] ),
    .Y(_12630_));
 sky130_fd_sc_hd__nand3_1 _17032_ (.A(_12586_),
    .B(_12588_),
    .C(_12601_),
    .Y(_12631_));
 sky130_fd_sc_hd__a21oi_1 _17033_ (.A1(_12603_),
    .A2(_12631_),
    .B1(\base_h_counter[3] ),
    .Y(_12632_));
 sky130_fd_sc_hd__nand3_1 _17034_ (.A(_12538_),
    .B(_12592_),
    .C(_12599_),
    .Y(_12633_));
 sky130_fd_sc_hd__a21oi_1 _17035_ (.A1(_12601_),
    .A2(_12633_),
    .B1(\base_h_counter[2] ),
    .Y(_12634_));
 sky130_fd_sc_hd__nand3_1 _17036_ (.A(_12601_),
    .B(_12633_),
    .C(\base_h_counter[2] ),
    .Y(_12635_));
 sky130_fd_sc_hd__nand3_1 _17037_ (.A(_12595_),
    .B(_12533_),
    .C(_12598_),
    .Y(_12636_));
 sky130_fd_sc_hd__nand3_1 _17038_ (.A(_12594_),
    .B(_12531_),
    .C(_12597_),
    .Y(_12637_));
 sky130_fd_sc_hd__nand2_1 _17039_ (.A(_12636_),
    .B(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand2_1 _17040_ (.A(_12638_),
    .B(\base_h_counter[1] ),
    .Y(_12639_));
 sky130_fd_sc_hd__xor2_1 _17041_ (.A(_08890_),
    .B(_12598_),
    .X(_12640_));
 sky130_fd_sc_hd__nand3_1 _17042_ (.A(_12636_),
    .B(_08891_),
    .C(_12637_),
    .Y(_12641_));
 sky130_fd_sc_hd__nand3_1 _17043_ (.A(_12639_),
    .B(_12640_),
    .C(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__inv_2 _17044_ (.A(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__nand2_1 _17045_ (.A(_12635_),
    .B(_12643_),
    .Y(_12644_));
 sky130_fd_sc_hd__nor2_1 _17046_ (.A(_12634_),
    .B(_12644_),
    .Y(_12645_));
 sky130_fd_sc_hd__nand3_1 _17047_ (.A(_12603_),
    .B(_12631_),
    .C(\base_h_counter[3] ),
    .Y(_12646_));
 sky130_fd_sc_hd__nand2_1 _17048_ (.A(_12645_),
    .B(_12646_),
    .Y(_12647_));
 sky130_fd_sc_hd__nor2_1 _17049_ (.A(_12632_),
    .B(_12647_),
    .Y(_12648_));
 sky130_fd_sc_hd__nand3_1 _17050_ (.A(_12605_),
    .B(_12629_),
    .C(\base_h_counter[4] ),
    .Y(_12649_));
 sky130_fd_sc_hd__nand2_1 _17051_ (.A(_12648_),
    .B(_12649_),
    .Y(_12650_));
 sky130_fd_sc_hd__nor2_1 _17052_ (.A(_12630_),
    .B(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__nand3_1 _17053_ (.A(_12605_),
    .B(_12579_),
    .C(_12572_),
    .Y(_12652_));
 sky130_fd_sc_hd__nand2_1 _17054_ (.A(_12607_),
    .B(_12652_),
    .Y(_12653_));
 sky130_fd_sc_hd__nand2_1 _17055_ (.A(_12653_),
    .B(_08885_),
    .Y(_12654_));
 sky130_fd_sc_hd__nand3_1 _17056_ (.A(_12607_),
    .B(_12652_),
    .C(\base_h_counter[5] ),
    .Y(_12655_));
 sky130_fd_sc_hd__nand3_1 _17057_ (.A(_12651_),
    .B(_12654_),
    .C(_12655_),
    .Y(_12656_));
 sky130_fd_sc_hd__nand3_1 _17058_ (.A(_12607_),
    .B(_12575_),
    .C(_12576_),
    .Y(_12657_));
 sky130_fd_sc_hd__nand2_1 _17059_ (.A(_12609_),
    .B(_12657_),
    .Y(_12658_));
 sky130_fd_sc_hd__nor2_1 _17060_ (.A(_08871_),
    .B(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__nor2_1 _17061_ (.A(_12656_),
    .B(_12659_),
    .Y(_12660_));
 sky130_fd_sc_hd__nand2_1 _17062_ (.A(_12658_),
    .B(_08871_),
    .Y(_12661_));
 sky130_fd_sc_hd__nand3_1 _17063_ (.A(_12628_),
    .B(_12660_),
    .C(_12661_),
    .Y(_12662_));
 sky130_fd_sc_hd__nor2_1 _17064_ (.A(_12627_),
    .B(_12662_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand2_1 _17065_ (.A(_12614_),
    .B(_12617_),
    .Y(_12664_));
 sky130_fd_sc_hd__inv_2 _17066_ (.A(_12617_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand2_1 _17067_ (.A(_12623_),
    .B(_12619_),
    .Y(_12666_));
 sky130_fd_sc_hd__nand2_1 _17068_ (.A(_12665_),
    .B(_12666_),
    .Y(_12667_));
 sky130_fd_sc_hd__nand3_1 _17069_ (.A(_12664_),
    .B(_12667_),
    .C(net3959),
    .Y(_12668_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(_12614_),
    .B(_12665_),
    .Y(_12669_));
 sky130_fd_sc_hd__nand2_1 _17071_ (.A(_12666_),
    .B(_12617_),
    .Y(_12670_));
 sky130_fd_sc_hd__nand3_1 _17072_ (.A(_12669_),
    .B(_08910_),
    .C(_12670_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand2_1 _17073_ (.A(_12668_),
    .B(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__inv_2 _17074_ (.A(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__inv_2 _17075_ (.A(_12566_),
    .Y(_12674_));
 sky130_fd_sc_hd__nand2_1 _17076_ (.A(_12664_),
    .B(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__nand2_1 _17077_ (.A(_12675_),
    .B(_09252_),
    .Y(_12676_));
 sky130_fd_sc_hd__nand3_1 _17078_ (.A(_12664_),
    .B(_12674_),
    .C(net3947),
    .Y(_12677_));
 sky130_fd_sc_hd__nand2_1 _17079_ (.A(_12676_),
    .B(_12677_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3_4 _17080_ (.A(_12663_),
    .B(_12673_),
    .C(_12678_),
    .Y(_12679_));
 sky130_fd_sc_hd__nand3_4 _17081_ (.A(_12679_),
    .B(_09126_),
    .C(_09114_),
    .Y(_12680_));
 sky130_fd_sc_hd__nand2_1 _17082_ (.A(_09498_),
    .B(net1985),
    .Y(_12681_));
 sky130_fd_sc_hd__o21ai_1 _17083_ (.A1(net1985),
    .A2(_12680_),
    .B1(_12681_),
    .Y(_00131_));
 sky130_fd_sc_hd__clkbuf_8 _17084_ (.A(_09496_),
    .X(_12682_));
 sky130_fd_sc_hd__nand2_1 _17085_ (.A(_08891_),
    .B(_08890_),
    .Y(_12683_));
 sky130_fd_sc_hd__nand2_2 _17086_ (.A(net3965),
    .B(net1985),
    .Y(_12684_));
 sky130_fd_sc_hd__nand2_1 _17087_ (.A(_12683_),
    .B(_12684_),
    .Y(_12685_));
 sky130_fd_sc_hd__buf_6 _17088_ (.A(_12680_),
    .X(_12686_));
 sky130_fd_sc_hd__o22ai_1 _17089_ (.A1(_08891_),
    .A2(_12682_),
    .B1(_12685_),
    .B2(_12686_),
    .Y(_00132_));
 sky130_fd_sc_hd__xor2_1 _17090_ (.A(net3976),
    .B(_12684_),
    .X(_12687_));
 sky130_fd_sc_hd__o22ai_1 _17091_ (.A1(_08898_),
    .A2(_12682_),
    .B1(_12687_),
    .B2(_12686_),
    .Y(_00133_));
 sky130_fd_sc_hd__nor3_1 _17092_ (.A(_08901_),
    .B(_08898_),
    .C(_12684_),
    .Y(_12688_));
 sky130_fd_sc_hd__o21ai_1 _17093_ (.A1(_08898_),
    .A2(_12684_),
    .B1(_08901_),
    .Y(_12689_));
 sky130_fd_sc_hd__or2b_1 _17094_ (.A(_12688_),
    .B_N(_12689_),
    .X(_12690_));
 sky130_fd_sc_hd__o22ai_1 _17095_ (.A1(_08901_),
    .A2(_12682_),
    .B1(_12690_),
    .B2(_12686_),
    .Y(_00134_));
 sky130_fd_sc_hd__or2_1 _17096_ (.A(net3994),
    .B(_12688_),
    .X(_12691_));
 sky130_fd_sc_hd__nand2_1 _17097_ (.A(_12688_),
    .B(net3994),
    .Y(_12692_));
 sky130_fd_sc_hd__nand2_1 _17098_ (.A(_12691_),
    .B(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__o22ai_1 _17099_ (.A1(_08879_),
    .A2(_09497_),
    .B1(_12693_),
    .B2(_12686_),
    .Y(_00135_));
 sky130_fd_sc_hd__or2_1 _17100_ (.A(_08885_),
    .B(_12692_),
    .X(_12694_));
 sky130_fd_sc_hd__nand2_1 _17101_ (.A(_12692_),
    .B(_08885_),
    .Y(_12695_));
 sky130_fd_sc_hd__nand2_1 _17102_ (.A(_12694_),
    .B(_12695_),
    .Y(_12696_));
 sky130_fd_sc_hd__o22ai_1 _17103_ (.A1(_08885_),
    .A2(_09497_),
    .B1(_12696_),
    .B2(_12686_),
    .Y(_00136_));
 sky130_fd_sc_hd__or2_1 _17104_ (.A(_08871_),
    .B(_12694_),
    .X(_12697_));
 sky130_fd_sc_hd__nand2_1 _17105_ (.A(_12694_),
    .B(_08871_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand2_1 _17106_ (.A(_12697_),
    .B(_12698_),
    .Y(_12699_));
 sky130_fd_sc_hd__o22ai_1 _17107_ (.A1(_08871_),
    .A2(_09497_),
    .B1(_12699_),
    .B2(_12686_),
    .Y(_00137_));
 sky130_fd_sc_hd__nor2_1 _17108_ (.A(_08874_),
    .B(_12697_),
    .Y(_12700_));
 sky130_fd_sc_hd__inv_2 _17109_ (.A(_12700_),
    .Y(_12701_));
 sky130_fd_sc_hd__nand2_1 _17110_ (.A(_12697_),
    .B(_08874_),
    .Y(_12702_));
 sky130_fd_sc_hd__nand2_1 _17111_ (.A(_12701_),
    .B(_12702_),
    .Y(_12703_));
 sky130_fd_sc_hd__o22ai_1 _17112_ (.A1(_08874_),
    .A2(_09497_),
    .B1(_12703_),
    .B2(_12680_),
    .Y(_00138_));
 sky130_fd_sc_hd__nor2_1 _17113_ (.A(net3959),
    .B(_12700_),
    .Y(_12704_));
 sky130_fd_sc_hd__nor2_1 _17114_ (.A(_08910_),
    .B(_12701_),
    .Y(_12705_));
 sky130_fd_sc_hd__or2_1 _17115_ (.A(_12704_),
    .B(_12705_),
    .X(_12706_));
 sky130_fd_sc_hd__o22ai_1 _17116_ (.A1(_08910_),
    .A2(_09497_),
    .B1(_12706_),
    .B2(_12680_),
    .Y(_00139_));
 sky130_fd_sc_hd__xor2_1 _17117_ (.A(_09252_),
    .B(_12705_),
    .X(_12707_));
 sky130_fd_sc_hd__o22ai_1 _17118_ (.A1(_09252_),
    .A2(_09497_),
    .B1(_12707_),
    .B2(_12680_),
    .Y(_00140_));
 sky130_fd_sc_hd__inv_2 _17119_ (.A(\base_v_bporch[2] ),
    .Y(_12708_));
 sky130_fd_sc_hd__nand2_1 _17120_ (.A(_09475_),
    .B(_12708_),
    .Y(_12709_));
 sky130_fd_sc_hd__nand3_2 _17121_ (.A(_09474_),
    .B(\base_v_bporch[2] ),
    .C(_09423_),
    .Y(_12710_));
 sky130_fd_sc_hd__nand2_1 _17122_ (.A(_09464_),
    .B(\base_v_bporch[0] ),
    .Y(_12711_));
 sky130_fd_sc_hd__inv_2 _17123_ (.A(\base_v_bporch[1] ),
    .Y(_12712_));
 sky130_fd_sc_hd__nand2_1 _17124_ (.A(_09467_),
    .B(_12712_),
    .Y(_12713_));
 sky130_fd_sc_hd__nand3_1 _17125_ (.A(_09466_),
    .B(\base_v_bporch[1] ),
    .C(_09418_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand3b_1 _17126_ (.A_N(_12711_),
    .B(_12713_),
    .C(_12714_),
    .Y(_12715_));
 sky130_fd_sc_hd__nand2_1 _17127_ (.A(_12715_),
    .B(_12714_),
    .Y(_12716_));
 sky130_fd_sc_hd__nand3_2 _17128_ (.A(_12709_),
    .B(_12710_),
    .C(_12716_),
    .Y(_12717_));
 sky130_fd_sc_hd__nand2_1 _17129_ (.A(_12717_),
    .B(_12710_),
    .Y(_12718_));
 sky130_fd_sc_hd__nand2b_2 _17130_ (.A_N(_09472_),
    .B(\base_v_bporch[3] ),
    .Y(_12719_));
 sky130_fd_sc_hd__a21o_1 _17131_ (.A1(_09425_),
    .A2(_09471_),
    .B1(\base_v_bporch[3] ),
    .X(_12720_));
 sky130_fd_sc_hd__nand3_2 _17132_ (.A(_12718_),
    .B(_12719_),
    .C(_12720_),
    .Y(_12721_));
 sky130_fd_sc_hd__nand2_1 _17133_ (.A(_12721_),
    .B(_12719_),
    .Y(_12722_));
 sky130_fd_sc_hd__nand2_1 _17134_ (.A(_12722_),
    .B(_09429_),
    .Y(_12723_));
 sky130_fd_sc_hd__nand3_1 _17135_ (.A(_12721_),
    .B(_09428_),
    .C(_12719_),
    .Y(_12724_));
 sky130_fd_sc_hd__nand2_1 _17136_ (.A(_12719_),
    .B(_12720_),
    .Y(_12725_));
 sky130_fd_sc_hd__nand3_1 _17137_ (.A(_12725_),
    .B(_12717_),
    .C(_12710_),
    .Y(_12726_));
 sky130_fd_sc_hd__nand2_1 _17138_ (.A(_12726_),
    .B(_12721_),
    .Y(_12727_));
 sky130_fd_sc_hd__nand2_1 _17139_ (.A(_12709_),
    .B(_12710_),
    .Y(_12728_));
 sky130_fd_sc_hd__inv_2 _17140_ (.A(_12716_),
    .Y(_12729_));
 sky130_fd_sc_hd__nand2_1 _17141_ (.A(_12728_),
    .B(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_1 _17142_ (.A(_12730_),
    .B(_12717_),
    .Y(_12731_));
 sky130_fd_sc_hd__nand2_1 _17143_ (.A(_12713_),
    .B(_12714_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand2_1 _17144_ (.A(_12732_),
    .B(_12711_),
    .Y(_12733_));
 sky130_fd_sc_hd__nand2_1 _17145_ (.A(_12733_),
    .B(_12715_),
    .Y(_12734_));
 sky130_fd_sc_hd__or2_1 _17146_ (.A(\base_v_bporch[0] ),
    .B(_09464_),
    .X(_12735_));
 sky130_fd_sc_hd__nand2_1 _17147_ (.A(_12735_),
    .B(_12711_),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(_12734_),
    .B(_12736_),
    .Y(_12737_));
 sky130_fd_sc_hd__inv_2 _17149_ (.A(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_1 _17150_ (.A(_12731_),
    .B(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__inv_2 _17151_ (.A(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_2 _17152_ (.A(_12727_),
    .B(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__a21oi_2 _17153_ (.A1(_12723_),
    .A2(_12724_),
    .B1(_12741_),
    .Y(_12742_));
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(_12723_),
    .B(_09435_),
    .Y(_12743_));
 sky130_fd_sc_hd__nand3_1 _17155_ (.A(_09426_),
    .B(_09370_),
    .C(_09427_),
    .Y(_12744_));
 sky130_fd_sc_hd__inv_2 _17156_ (.A(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__nand2_1 _17157_ (.A(_12722_),
    .B(_12745_),
    .Y(_12746_));
 sky130_fd_sc_hd__nand2_2 _17158_ (.A(_12743_),
    .B(_12746_),
    .Y(_12747_));
 sky130_fd_sc_hd__nand2_1 _17159_ (.A(_12746_),
    .B(_09447_),
    .Y(_12748_));
 sky130_fd_sc_hd__nand3b_1 _17160_ (.A_N(_09447_),
    .B(_12722_),
    .C(_12745_),
    .Y(_12749_));
 sky130_fd_sc_hd__nand2_1 _17161_ (.A(_12748_),
    .B(_12749_),
    .Y(_12750_));
 sky130_fd_sc_hd__nand3_2 _17162_ (.A(_12742_),
    .B(_12747_),
    .C(_12750_),
    .Y(_12751_));
 sky130_fd_sc_hd__inv_2 _17163_ (.A(_12751_),
    .Y(_12752_));
 sky130_fd_sc_hd__nand2_1 _17164_ (.A(_12749_),
    .B(_09444_),
    .Y(_12753_));
 sky130_fd_sc_hd__nand3_1 _17165_ (.A(_09441_),
    .B(_09403_),
    .C(_09446_),
    .Y(_12754_));
 sky130_fd_sc_hd__nand3b_1 _17166_ (.A_N(_12754_),
    .B(_12722_),
    .C(_12745_),
    .Y(_12755_));
 sky130_fd_sc_hd__nand2_1 _17167_ (.A(_12753_),
    .B(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__nand2_1 _17168_ (.A(_12752_),
    .B(_12756_),
    .Y(_12757_));
 sky130_fd_sc_hd__inv_2 _17169_ (.A(_12756_),
    .Y(_12758_));
 sky130_fd_sc_hd__nand2_1 _17170_ (.A(_12751_),
    .B(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(_12757_),
    .B(_12759_),
    .Y(_12760_));
 sky130_fd_sc_hd__nand2_1 _17172_ (.A(_12760_),
    .B(_08920_),
    .Y(_12761_));
 sky130_fd_sc_hd__nand3_1 _17173_ (.A(_12757_),
    .B(_08919_),
    .C(_12759_),
    .Y(_12762_));
 sky130_fd_sc_hd__or2_1 _17174_ (.A(_09457_),
    .B(_12755_),
    .X(_12763_));
 sky130_fd_sc_hd__nand2_1 _17175_ (.A(_12763_),
    .B(_09491_),
    .Y(_12764_));
 sky130_fd_sc_hd__or2_1 _17176_ (.A(_08960_),
    .B(_12764_),
    .X(_12765_));
 sky130_fd_sc_hd__nand3_1 _17177_ (.A(_12761_),
    .B(_12762_),
    .C(_12765_),
    .Y(_12766_));
 sky130_fd_sc_hd__nand2_1 _17178_ (.A(_12742_),
    .B(_12747_),
    .Y(_12767_));
 sky130_fd_sc_hd__inv_2 _17179_ (.A(_12750_),
    .Y(_12768_));
 sky130_fd_sc_hd__nand2_1 _17180_ (.A(_12767_),
    .B(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(_12769_),
    .B(_12751_),
    .Y(_12770_));
 sky130_fd_sc_hd__nand2_1 _17182_ (.A(_12770_),
    .B(_08917_),
    .Y(_12771_));
 sky130_fd_sc_hd__nand3_1 _17183_ (.A(_12769_),
    .B(net3812),
    .C(_12751_),
    .Y(_12772_));
 sky130_fd_sc_hd__nand2_1 _17184_ (.A(_12771_),
    .B(_12772_),
    .Y(_12773_));
 sky130_fd_sc_hd__inv_2 _17185_ (.A(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__nand3_1 _17186_ (.A(_12726_),
    .B(_12721_),
    .C(_12739_),
    .Y(_12775_));
 sky130_fd_sc_hd__a21oi_1 _17187_ (.A1(_12741_),
    .A2(_12775_),
    .B1(\base_v_counter[3] ),
    .Y(_12776_));
 sky130_fd_sc_hd__nand3_1 _17188_ (.A(_12730_),
    .B(_12717_),
    .C(_12737_),
    .Y(_12777_));
 sky130_fd_sc_hd__nand2_1 _17189_ (.A(_12739_),
    .B(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__and2_1 _17190_ (.A(_12778_),
    .B(_08949_),
    .X(_12779_));
 sky130_fd_sc_hd__or2b_1 _17191_ (.A(_12734_),
    .B_N(_12736_),
    .X(_12780_));
 sky130_fd_sc_hd__or2b_1 _17192_ (.A(_12736_),
    .B_N(_12734_),
    .X(_12781_));
 sky130_fd_sc_hd__nand2_1 _17193_ (.A(_12780_),
    .B(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__nand2_1 _17194_ (.A(_12782_),
    .B(\base_v_counter[1] ),
    .Y(_12783_));
 sky130_fd_sc_hd__nand3_1 _17195_ (.A(_12780_),
    .B(_12781_),
    .C(_09340_),
    .Y(_12784_));
 sky130_fd_sc_hd__xor2_1 _17196_ (.A(_08938_),
    .B(_12736_),
    .X(_12785_));
 sky130_fd_sc_hd__nand3_1 _17197_ (.A(_12783_),
    .B(_12784_),
    .C(_12785_),
    .Y(_12786_));
 sky130_fd_sc_hd__inv_2 _17198_ (.A(_12786_),
    .Y(_12787_));
 sky130_fd_sc_hd__o21ai_1 _17199_ (.A1(_08949_),
    .A2(_12778_),
    .B1(_12787_),
    .Y(_12788_));
 sky130_fd_sc_hd__nor2_1 _17200_ (.A(_12779_),
    .B(_12788_),
    .Y(_12789_));
 sky130_fd_sc_hd__nand3_1 _17201_ (.A(_12741_),
    .B(_12775_),
    .C(\base_v_counter[3] ),
    .Y(_12790_));
 sky130_fd_sc_hd__nand2_1 _17202_ (.A(_12789_),
    .B(_12790_),
    .Y(_12791_));
 sky130_fd_sc_hd__nor2_1 _17203_ (.A(_12776_),
    .B(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__nand2_1 _17204_ (.A(_12723_),
    .B(_12724_),
    .Y(_12793_));
 sky130_fd_sc_hd__inv_2 _17205_ (.A(_12793_),
    .Y(_12794_));
 sky130_fd_sc_hd__nand2_1 _17206_ (.A(_12794_),
    .B(_12741_),
    .Y(_12795_));
 sky130_fd_sc_hd__inv_2 _17207_ (.A(_12741_),
    .Y(_12796_));
 sky130_fd_sc_hd__nand2_1 _17208_ (.A(_12796_),
    .B(_12793_),
    .Y(_12797_));
 sky130_fd_sc_hd__nand2_1 _17209_ (.A(_12795_),
    .B(_12797_),
    .Y(_12798_));
 sky130_fd_sc_hd__nand2_1 _17210_ (.A(_12798_),
    .B(_08934_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand3_1 _17211_ (.A(_12795_),
    .B(net3797),
    .C(_12797_),
    .Y(_12800_));
 sky130_fd_sc_hd__nand3_1 _17212_ (.A(_12792_),
    .B(_12799_),
    .C(_12800_),
    .Y(_12801_));
 sky130_fd_sc_hd__inv_2 _17213_ (.A(_12747_),
    .Y(_12802_));
 sky130_fd_sc_hd__nand2_1 _17214_ (.A(_12802_),
    .B(_12742_),
    .Y(_12803_));
 sky130_fd_sc_hd__nand2_1 _17215_ (.A(_12797_),
    .B(_12747_),
    .Y(_12804_));
 sky130_fd_sc_hd__nand2_1 _17216_ (.A(_12803_),
    .B(_12804_),
    .Y(_12805_));
 sky130_fd_sc_hd__nand2_1 _17217_ (.A(_12805_),
    .B(net3817),
    .Y(_12806_));
 sky130_fd_sc_hd__nand3_1 _17218_ (.A(_12803_),
    .B(_08929_),
    .C(_12804_),
    .Y(_12807_));
 sky130_fd_sc_hd__nand2_1 _17219_ (.A(_12806_),
    .B(_12807_),
    .Y(_12808_));
 sky130_fd_sc_hd__nor2_1 _17220_ (.A(_12801_),
    .B(_12808_),
    .Y(_12809_));
 sky130_fd_sc_hd__nand2_1 _17221_ (.A(_12764_),
    .B(_08960_),
    .Y(_12810_));
 sky130_fd_sc_hd__nor2_1 _17222_ (.A(_12758_),
    .B(_12751_),
    .Y(_12811_));
 sky130_fd_sc_hd__nand2_1 _17223_ (.A(_12755_),
    .B(_09457_),
    .Y(_12812_));
 sky130_fd_sc_hd__nand2_1 _17224_ (.A(_12763_),
    .B(_12812_),
    .Y(_12813_));
 sky130_fd_sc_hd__nand3_1 _17225_ (.A(_12810_),
    .B(_12811_),
    .C(_12813_),
    .Y(_12814_));
 sky130_fd_sc_hd__nand3_1 _17226_ (.A(_12774_),
    .B(_12809_),
    .C(_12814_),
    .Y(_12815_));
 sky130_fd_sc_hd__nor2_1 _17227_ (.A(_12766_),
    .B(_12815_),
    .Y(_12816_));
 sky130_fd_sc_hd__inv_2 _17228_ (.A(_12813_),
    .Y(_12817_));
 sky130_fd_sc_hd__nand2_1 _17229_ (.A(_12757_),
    .B(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__nand2_1 _17230_ (.A(_12811_),
    .B(_12813_),
    .Y(_12819_));
 sky130_fd_sc_hd__a21oi_1 _17231_ (.A1(_12818_),
    .A2(_12819_),
    .B1(net3823),
    .Y(_12820_));
 sky130_fd_sc_hd__nand2b_1 _17232_ (.A_N(_12810_),
    .B(_12819_),
    .Y(_12821_));
 sky130_fd_sc_hd__nand3_1 _17233_ (.A(_12818_),
    .B(_12819_),
    .C(net3823),
    .Y(_12822_));
 sky130_fd_sc_hd__nand2_1 _17234_ (.A(_12821_),
    .B(_12822_),
    .Y(_12823_));
 sky130_fd_sc_hd__nor2_1 _17235_ (.A(_12820_),
    .B(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__nand2_4 _17236_ (.A(_12816_),
    .B(_12824_),
    .Y(_12825_));
 sky130_fd_sc_hd__nor2_1 _17237_ (.A(net2025),
    .B(_09130_),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2_1 _17238_ (.A(_12825_),
    .B(_12826_),
    .Y(_12827_));
 sky130_fd_sc_hd__or2_1 _17239_ (.A(net43),
    .B(net30),
    .X(_12828_));
 sky130_fd_sc_hd__nand2_1 _17240_ (.A(net43),
    .B(net30),
    .Y(_12829_));
 sky130_fd_sc_hd__nand2_1 _17241_ (.A(_12828_),
    .B(_12829_),
    .Y(_12830_));
 sky130_fd_sc_hd__inv_2 _17242_ (.A(_12830_),
    .Y(_12831_));
 sky130_fd_sc_hd__nor2_1 _17243_ (.A(net46),
    .B(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__nand2_1 _17244_ (.A(_12831_),
    .B(net46),
    .Y(_12833_));
 sky130_fd_sc_hd__or3b_1 _17245_ (.A(_09126_),
    .B(_12832_),
    .C_N(_12833_),
    .X(_12834_));
 sky130_fd_sc_hd__nand2_1 _17246_ (.A(_12827_),
    .B(_12834_),
    .Y(_12835_));
 sky130_fd_sc_hd__nand3_1 _17247_ (.A(_12835_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12836_));
 sky130_fd_sc_hd__nand2_4 _17248_ (.A(_12680_),
    .B(_09497_),
    .Y(_12837_));
 sky130_fd_sc_hd__nand2_1 _17249_ (.A(_12837_),
    .B(net2025),
    .Y(_12838_));
 sky130_fd_sc_hd__nand2_1 _17250_ (.A(_12836_),
    .B(net2026),
    .Y(_00141_));
 sky130_fd_sc_hd__nand2_1 _17251_ (.A(_09340_),
    .B(_08938_),
    .Y(_12839_));
 sky130_fd_sc_hd__clkbuf_8 _17252_ (.A(_09125_),
    .X(_12840_));
 sky130_fd_sc_hd__nand2_1 _17253_ (.A(net3800),
    .B(net2025),
    .Y(_12841_));
 sky130_fd_sc_hd__and3_1 _17254_ (.A(_12839_),
    .B(_12840_),
    .C(_12841_),
    .X(_12842_));
 sky130_fd_sc_hd__nand2_1 _17255_ (.A(_12825_),
    .B(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__and2_1 _17256_ (.A(_12833_),
    .B(_12829_),
    .X(_12844_));
 sky130_fd_sc_hd__or2_1 _17257_ (.A(net44),
    .B(net31),
    .X(_12845_));
 sky130_fd_sc_hd__nand2_1 _17258_ (.A(net44),
    .B(net31),
    .Y(_12846_));
 sky130_fd_sc_hd__nand2_1 _17259_ (.A(_12845_),
    .B(_12846_),
    .Y(_12847_));
 sky130_fd_sc_hd__xor2_1 _17260_ (.A(net47),
    .B(_12847_),
    .X(_12848_));
 sky130_fd_sc_hd__nor2_1 _17261_ (.A(_12848_),
    .B(_12844_),
    .Y(_12849_));
 sky130_fd_sc_hd__inv_2 _17262_ (.A(_12849_),
    .Y(_12850_));
 sky130_fd_sc_hd__buf_8 _17263_ (.A(_09057_),
    .X(_12851_));
 sky130_fd_sc_hd__nand2_1 _17264_ (.A(_12850_),
    .B(_12851_),
    .Y(_12852_));
 sky130_fd_sc_hd__a21o_1 _17265_ (.A1(_12844_),
    .A2(_12848_),
    .B1(_12852_),
    .X(_12853_));
 sky130_fd_sc_hd__nand2_1 _17266_ (.A(_12843_),
    .B(_12853_),
    .Y(_12854_));
 sky130_fd_sc_hd__nand3_1 _17267_ (.A(_12854_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12855_));
 sky130_fd_sc_hd__nand2_1 _17268_ (.A(_12837_),
    .B(net3800),
    .Y(_12856_));
 sky130_fd_sc_hd__nand2_1 _17269_ (.A(_12855_),
    .B(net3801),
    .Y(_00142_));
 sky130_fd_sc_hd__nor2_1 _17270_ (.A(_08949_),
    .B(_12841_),
    .Y(_12857_));
 sky130_fd_sc_hd__inv_2 _17271_ (.A(_12857_),
    .Y(_12858_));
 sky130_fd_sc_hd__nand2_1 _17272_ (.A(_12841_),
    .B(_08949_),
    .Y(_12859_));
 sky130_fd_sc_hd__and3_1 _17273_ (.A(_12858_),
    .B(_12840_),
    .C(_12859_),
    .X(_12860_));
 sky130_fd_sc_hd__nand2_1 _17274_ (.A(_12825_),
    .B(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__a21boi_1 _17275_ (.A1(_12845_),
    .A2(net47),
    .B1_N(_12846_),
    .Y(_12862_));
 sky130_fd_sc_hd__inv_2 _17276_ (.A(net48),
    .Y(_12863_));
 sky130_fd_sc_hd__or2_1 _17277_ (.A(net45),
    .B(net32),
    .X(_12864_));
 sky130_fd_sc_hd__nand2_1 _17278_ (.A(net45),
    .B(net32),
    .Y(_12865_));
 sky130_fd_sc_hd__nand2_1 _17279_ (.A(_12864_),
    .B(_12865_),
    .Y(_12866_));
 sky130_fd_sc_hd__or2_1 _17280_ (.A(_12863_),
    .B(_12866_),
    .X(_12867_));
 sky130_fd_sc_hd__nand2_1 _17281_ (.A(_12866_),
    .B(_12863_),
    .Y(_12868_));
 sky130_fd_sc_hd__nand2_1 _17282_ (.A(_12867_),
    .B(_12868_),
    .Y(_12869_));
 sky130_fd_sc_hd__or2_1 _17283_ (.A(_12862_),
    .B(_12869_),
    .X(_12870_));
 sky130_fd_sc_hd__nand2_1 _17284_ (.A(_12869_),
    .B(_12862_),
    .Y(_12871_));
 sky130_fd_sc_hd__nand2_1 _17285_ (.A(_12870_),
    .B(_12871_),
    .Y(_12872_));
 sky130_fd_sc_hd__or2_1 _17286_ (.A(_12850_),
    .B(_12872_),
    .X(_12873_));
 sky130_fd_sc_hd__nand2_1 _17287_ (.A(_12873_),
    .B(_12851_),
    .Y(_12874_));
 sky130_fd_sc_hd__a21o_1 _17288_ (.A1(_12850_),
    .A2(_12872_),
    .B1(_12874_),
    .X(_12875_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(_12861_),
    .B(_12875_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand3_1 _17290_ (.A(_12876_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12877_));
 sky130_fd_sc_hd__nand2_1 _17291_ (.A(_12837_),
    .B(net2011),
    .Y(_12878_));
 sky130_fd_sc_hd__nand2_1 _17292_ (.A(_12877_),
    .B(net2012),
    .Y(_00143_));
 sky130_fd_sc_hd__nor2_1 _17293_ (.A(_08944_),
    .B(_12858_),
    .Y(_12879_));
 sky130_fd_sc_hd__inv_2 _17294_ (.A(_12879_),
    .Y(_12880_));
 sky130_fd_sc_hd__nand2_1 _17295_ (.A(_12858_),
    .B(_08944_),
    .Y(_12881_));
 sky130_fd_sc_hd__and3_1 _17296_ (.A(_12880_),
    .B(_12840_),
    .C(_12881_),
    .X(_12882_));
 sky130_fd_sc_hd__nand2_1 _17297_ (.A(_12825_),
    .B(_12882_),
    .Y(_12883_));
 sky130_fd_sc_hd__nand2_1 _17298_ (.A(_12867_),
    .B(_12865_),
    .Y(_12884_));
 sky130_fd_sc_hd__inv_2 _17299_ (.A(_12884_),
    .Y(_12885_));
 sky130_fd_sc_hd__nor2_1 _17300_ (.A(_12269_),
    .B(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__nand2_1 _17301_ (.A(_12885_),
    .B(_12269_),
    .Y(_12887_));
 sky130_fd_sc_hd__or2b_1 _17302_ (.A(_12886_),
    .B_N(_12887_),
    .X(_12888_));
 sky130_fd_sc_hd__nand2_2 _17303_ (.A(_12873_),
    .B(_12870_),
    .Y(_12889_));
 sky130_fd_sc_hd__or2_1 _17304_ (.A(_12888_),
    .B(_12889_),
    .X(_12890_));
 sky130_fd_sc_hd__nand2_1 _17305_ (.A(_12889_),
    .B(_12888_),
    .Y(_12891_));
 sky130_fd_sc_hd__a21o_1 _17306_ (.A1(_12890_),
    .A2(_12891_),
    .B1(_09516_),
    .X(_12892_));
 sky130_fd_sc_hd__nand2_1 _17307_ (.A(_12883_),
    .B(_12892_),
    .Y(_12893_));
 sky130_fd_sc_hd__nand3_1 _17308_ (.A(_12893_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12894_));
 sky130_fd_sc_hd__nand2_1 _17309_ (.A(_12837_),
    .B(net3784),
    .Y(_12895_));
 sky130_fd_sc_hd__nand2_1 _17310_ (.A(_12894_),
    .B(net3785),
    .Y(_00144_));
 sky130_fd_sc_hd__nor2_1 _17311_ (.A(net3797),
    .B(_12879_),
    .Y(_12896_));
 sky130_fd_sc_hd__nor2_1 _17312_ (.A(_08934_),
    .B(_12880_),
    .Y(_12897_));
 sky130_fd_sc_hd__or3_1 _17313_ (.A(_09057_),
    .B(_12896_),
    .C(_12897_),
    .X(_12898_));
 sky130_fd_sc_hd__inv_2 _17314_ (.A(_12898_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand2_1 _17315_ (.A(_12825_),
    .B(_12899_),
    .Y(_12900_));
 sky130_fd_sc_hd__a21o_1 _17316_ (.A1(_12889_),
    .A2(_12887_),
    .B1(_12886_),
    .X(_12901_));
 sky130_fd_sc_hd__or2_1 _17317_ (.A(net34),
    .B(_12901_),
    .X(_12902_));
 sky130_fd_sc_hd__nand2_1 _17318_ (.A(_12901_),
    .B(net34),
    .Y(_12903_));
 sky130_fd_sc_hd__nand3_1 _17319_ (.A(_12902_),
    .B(_09130_),
    .C(_12903_),
    .Y(_12904_));
 sky130_fd_sc_hd__nand2_1 _17320_ (.A(_12900_),
    .B(_12904_),
    .Y(_12905_));
 sky130_fd_sc_hd__nand3_1 _17321_ (.A(_12905_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12906_));
 sky130_fd_sc_hd__nand2_1 _17322_ (.A(_12837_),
    .B(net3797),
    .Y(_12907_));
 sky130_fd_sc_hd__nand2_1 _17323_ (.A(_12906_),
    .B(net3798),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _17324_ (.A(_12897_),
    .Y(_12908_));
 sky130_fd_sc_hd__nor2_1 _17325_ (.A(_08929_),
    .B(_12908_),
    .Y(_12909_));
 sky130_fd_sc_hd__nor2_1 _17326_ (.A(_12851_),
    .B(_12909_),
    .Y(_12910_));
 sky130_fd_sc_hd__o21a_1 _17327_ (.A1(net3817),
    .A2(_12897_),
    .B1(_12910_),
    .X(_12911_));
 sky130_fd_sc_hd__nand2_1 _17328_ (.A(_12825_),
    .B(_12911_),
    .Y(_12912_));
 sky130_fd_sc_hd__nor2_1 _17329_ (.A(_12276_),
    .B(_12903_),
    .Y(_12913_));
 sky130_fd_sc_hd__or2_1 _17330_ (.A(_09126_),
    .B(_12913_),
    .X(_12914_));
 sky130_fd_sc_hd__a21o_1 _17331_ (.A1(_12276_),
    .A2(_12903_),
    .B1(_12914_),
    .X(_12915_));
 sky130_fd_sc_hd__nand2_1 _17332_ (.A(_12912_),
    .B(_12915_),
    .Y(_12916_));
 sky130_fd_sc_hd__nand3_1 _17333_ (.A(_12916_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12917_));
 sky130_fd_sc_hd__nand2_1 _17334_ (.A(_12837_),
    .B(net3817),
    .Y(_12918_));
 sky130_fd_sc_hd__nand2_1 _17335_ (.A(_12917_),
    .B(net3818),
    .Y(_00146_));
 sky130_fd_sc_hd__nor2_1 _17336_ (.A(net3812),
    .B(_12909_),
    .Y(_12919_));
 sky130_fd_sc_hd__nand2_1 _17337_ (.A(_12909_),
    .B(net3812),
    .Y(_12920_));
 sky130_fd_sc_hd__or3b_1 _17338_ (.A(_09057_),
    .B(_12919_),
    .C_N(_12920_),
    .X(_12921_));
 sky130_fd_sc_hd__inv_2 _17339_ (.A(_12921_),
    .Y(_12922_));
 sky130_fd_sc_hd__nand2_1 _17340_ (.A(_12825_),
    .B(_12922_),
    .Y(_12923_));
 sky130_fd_sc_hd__nor2_1 _17341_ (.A(net36),
    .B(_12913_),
    .Y(_12924_));
 sky130_fd_sc_hd__nand2_1 _17342_ (.A(_12913_),
    .B(net36),
    .Y(_12925_));
 sky130_fd_sc_hd__inv_2 _17343_ (.A(_12925_),
    .Y(_12926_));
 sky130_fd_sc_hd__or3_1 _17344_ (.A(_09126_),
    .B(_12924_),
    .C(_12926_),
    .X(_12927_));
 sky130_fd_sc_hd__nand2_1 _17345_ (.A(_12923_),
    .B(_12927_),
    .Y(_12928_));
 sky130_fd_sc_hd__nand3_1 _17346_ (.A(_12928_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12929_));
 sky130_fd_sc_hd__nand2_1 _17347_ (.A(_12837_),
    .B(net3812),
    .Y(_12930_));
 sky130_fd_sc_hd__nand2_1 _17348_ (.A(_12929_),
    .B(net3813),
    .Y(_00147_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(_08920_),
    .B(_12920_),
    .Y(_12931_));
 sky130_fd_sc_hd__nand2_1 _17350_ (.A(_12920_),
    .B(_08920_),
    .Y(_12932_));
 sky130_fd_sc_hd__or3b_1 _17351_ (.A(_09057_),
    .B(_12931_),
    .C_N(_12932_),
    .X(_12933_));
 sky130_fd_sc_hd__inv_2 _17352_ (.A(_12933_),
    .Y(_12934_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(_12825_),
    .B(_12934_),
    .Y(_12935_));
 sky130_fd_sc_hd__inv_2 _17354_ (.A(net37),
    .Y(_12936_));
 sky130_fd_sc_hd__nor2_1 _17355_ (.A(_12936_),
    .B(_12925_),
    .Y(_12937_));
 sky130_fd_sc_hd__nor2_1 _17356_ (.A(_09516_),
    .B(_12937_),
    .Y(_12938_));
 sky130_fd_sc_hd__o21ai_1 _17357_ (.A1(net37),
    .A2(_12926_),
    .B1(_12938_),
    .Y(_12939_));
 sky130_fd_sc_hd__nand2_1 _17358_ (.A(_12935_),
    .B(_12939_),
    .Y(_12940_));
 sky130_fd_sc_hd__nand3_1 _17359_ (.A(_12940_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12941_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(_12837_),
    .B(_08919_),
    .Y(_12942_));
 sky130_fd_sc_hd__nand2_1 _17361_ (.A(_12941_),
    .B(net3937),
    .Y(_00148_));
 sky130_fd_sc_hd__or2_1 _17362_ (.A(net3823),
    .B(_12931_),
    .X(_12943_));
 sky130_fd_sc_hd__nand2_1 _17363_ (.A(_12931_),
    .B(net3823),
    .Y(_12944_));
 sky130_fd_sc_hd__and3_1 _17364_ (.A(_12943_),
    .B(_12840_),
    .C(_12944_),
    .X(_12945_));
 sky130_fd_sc_hd__nand2_1 _17365_ (.A(_12825_),
    .B(_12945_),
    .Y(_12946_));
 sky130_fd_sc_hd__inv_2 _17366_ (.A(_12937_),
    .Y(_12947_));
 sky130_fd_sc_hd__a21o_1 _17367_ (.A1(_12937_),
    .A2(net38),
    .B1(_09126_),
    .X(_12948_));
 sky130_fd_sc_hd__a21o_1 _17368_ (.A1(_12285_),
    .A2(_12947_),
    .B1(_12948_),
    .X(_12949_));
 sky130_fd_sc_hd__nand2_1 _17369_ (.A(_12946_),
    .B(_12949_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand3_1 _17370_ (.A(_12950_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12951_));
 sky130_fd_sc_hd__nand2_1 _17371_ (.A(_12837_),
    .B(net3823),
    .Y(_12952_));
 sky130_fd_sc_hd__nand2_1 _17372_ (.A(_12951_),
    .B(net3824),
    .Y(_00149_));
 sky130_fd_sc_hd__a21oi_1 _17373_ (.A1(_12944_),
    .A2(_08960_),
    .B1(_12851_),
    .Y(_12953_));
 sky130_fd_sc_hd__o21a_1 _17374_ (.A1(_08960_),
    .A2(_12944_),
    .B1(_12953_),
    .X(_12954_));
 sky130_fd_sc_hd__nand2_1 _17375_ (.A(_12825_),
    .B(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__or3_1 _17376_ (.A(_09126_),
    .B(_12285_),
    .C(_12947_),
    .X(_12956_));
 sky130_fd_sc_hd__nand2_1 _17377_ (.A(_12955_),
    .B(_12956_),
    .Y(_12957_));
 sky130_fd_sc_hd__nand3_1 _17378_ (.A(_12957_),
    .B(_12686_),
    .C(_12682_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand2_1 _17379_ (.A(_12837_),
    .B(net3713),
    .Y(_12959_));
 sky130_fd_sc_hd__nand2_1 _17380_ (.A(_12958_),
    .B(net3714),
    .Y(_00150_));
 sky130_fd_sc_hd__buf_6 _17381_ (.A(_12679_),
    .X(_12960_));
 sky130_fd_sc_hd__nand2_1 _17382_ (.A(_09052_),
    .B(_09126_),
    .Y(_12961_));
 sky130_fd_sc_hd__inv_2 _17383_ (.A(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__nand3_1 _17384_ (.A(_12960_),
    .B(_09017_),
    .C(_12962_),
    .Y(_12963_));
 sky130_fd_sc_hd__nand2_1 _17385_ (.A(_08977_),
    .B(net49),
    .Y(_12964_));
 sky130_fd_sc_hd__inv_2 _17386_ (.A(_12964_),
    .Y(_12965_));
 sky130_fd_sc_hd__nand3_2 _17387_ (.A(_12679_),
    .B(_09114_),
    .C(_12965_),
    .Y(_12966_));
 sky130_fd_sc_hd__nor2_1 _17388_ (.A(_09056_),
    .B(_08869_),
    .Y(_12967_));
 sky130_fd_sc_hd__inv_2 _17389_ (.A(_12967_),
    .Y(_12968_));
 sky130_fd_sc_hd__nor2_1 _17390_ (.A(_12968_),
    .B(_09131_),
    .Y(_12969_));
 sky130_fd_sc_hd__nand2_1 _17391_ (.A(_12679_),
    .B(_12969_),
    .Y(_12970_));
 sky130_fd_sc_hd__nand3_4 _17392_ (.A(_12966_),
    .B(_09496_),
    .C(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__buf_6 _17393_ (.A(_12971_),
    .X(_12972_));
 sky130_fd_sc_hd__nand2_1 _17394_ (.A(_12972_),
    .B(net3773),
    .Y(_12973_));
 sky130_fd_sc_hd__o21ai_1 _17395_ (.A1(_12963_),
    .A2(_12972_),
    .B1(_12973_),
    .Y(_00151_));
 sky130_fd_sc_hd__o211ai_1 _17396_ (.A1(_09556_),
    .A2(_09566_),
    .B1(_12962_),
    .C1(_12960_),
    .Y(_12974_));
 sky130_fd_sc_hd__nand2_1 _17397_ (.A(_12972_),
    .B(net3867),
    .Y(_12975_));
 sky130_fd_sc_hd__o21ai_1 _17398_ (.A1(_12974_),
    .A2(_12972_),
    .B1(_12975_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_1 _17399_ (.A(_09562_),
    .B(net3745),
    .Y(_12976_));
 sky130_fd_sc_hd__nand2_1 _17400_ (.A(_09561_),
    .B(_09029_),
    .Y(_12977_));
 sky130_fd_sc_hd__and3_1 _17401_ (.A(_12976_),
    .B(_12840_),
    .C(_12977_),
    .X(_12978_));
 sky130_fd_sc_hd__nand3_1 _17402_ (.A(_12960_),
    .B(_09052_),
    .C(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__nand2_1 _17403_ (.A(_12972_),
    .B(net3745),
    .Y(_12980_));
 sky130_fd_sc_hd__o21ai_1 _17404_ (.A1(_12979_),
    .A2(_12972_),
    .B1(_12980_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_1 _17405_ (.A(_12976_),
    .B(_09021_),
    .Y(_12981_));
 sky130_fd_sc_hd__and3_1 _17406_ (.A(_12981_),
    .B(_12840_),
    .C(_09601_),
    .X(_12982_));
 sky130_fd_sc_hd__nand3_1 _17407_ (.A(_12960_),
    .B(_09052_),
    .C(_12982_),
    .Y(_12983_));
 sky130_fd_sc_hd__nand2_1 _17408_ (.A(_12972_),
    .B(net3638),
    .Y(_12984_));
 sky130_fd_sc_hd__o21ai_1 _17409_ (.A1(_12983_),
    .A2(_12972_),
    .B1(_12984_),
    .Y(_00154_));
 sky130_fd_sc_hd__nor2_1 _17410_ (.A(net3943),
    .B(_10109_),
    .Y(_12985_));
 sky130_fd_sc_hd__nor2_1 _17411_ (.A(_09047_),
    .B(_09601_),
    .Y(_12986_));
 sky130_fd_sc_hd__nor2_1 _17412_ (.A(_12985_),
    .B(_12986_),
    .Y(_12987_));
 sky130_fd_sc_hd__nand3_1 _17413_ (.A(_12960_),
    .B(_12962_),
    .C(_12987_),
    .Y(_12988_));
 sky130_fd_sc_hd__nand2_1 _17414_ (.A(_12972_),
    .B(net3943),
    .Y(_12989_));
 sky130_fd_sc_hd__o21ai_1 _17415_ (.A1(_12988_),
    .A2(_12972_),
    .B1(_12989_),
    .Y(_00155_));
 sky130_fd_sc_hd__or2_1 _17416_ (.A(net3902),
    .B(_12986_),
    .X(_12990_));
 sky130_fd_sc_hd__nand2_1 _17417_ (.A(_10109_),
    .B(_09553_),
    .Y(_12991_));
 sky130_fd_sc_hd__and3_1 _17418_ (.A(_12990_),
    .B(_12840_),
    .C(_12991_),
    .X(_12992_));
 sky130_fd_sc_hd__nand3_1 _17419_ (.A(_12960_),
    .B(_09052_),
    .C(_12992_),
    .Y(_12993_));
 sky130_fd_sc_hd__nand2_1 _17420_ (.A(_12972_),
    .B(net3902),
    .Y(_12994_));
 sky130_fd_sc_hd__o21ai_1 _17421_ (.A1(_12993_),
    .A2(_12972_),
    .B1(_12994_),
    .Y(_00156_));
 sky130_fd_sc_hd__or2_1 _17422_ (.A(_09013_),
    .B(_12991_),
    .X(_12995_));
 sky130_fd_sc_hd__nand2_1 _17423_ (.A(_12991_),
    .B(_09013_),
    .Y(_12996_));
 sky130_fd_sc_hd__and3_1 _17424_ (.A(_12995_),
    .B(_12840_),
    .C(_12996_),
    .X(_12997_));
 sky130_fd_sc_hd__nand3_1 _17425_ (.A(_12960_),
    .B(_09052_),
    .C(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__nand2_1 _17426_ (.A(_12972_),
    .B(net1997),
    .Y(_12999_));
 sky130_fd_sc_hd__o21ai_1 _17427_ (.A1(_12998_),
    .A2(_12971_),
    .B1(_12999_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _17428_ (.A(_12995_),
    .B(_09035_),
    .Y(_13000_));
 sky130_fd_sc_hd__and3_1 _17429_ (.A(_13000_),
    .B(_09126_),
    .C(_09603_),
    .X(_13001_));
 sky130_fd_sc_hd__nand3_1 _17430_ (.A(_12960_),
    .B(_09052_),
    .C(_13001_),
    .Y(_13002_));
 sky130_fd_sc_hd__nand2_1 _17431_ (.A(_12972_),
    .B(net3915),
    .Y(_13003_));
 sky130_fd_sc_hd__o21ai_1 _17432_ (.A1(_13002_),
    .A2(_12971_),
    .B1(_13003_),
    .Y(_00158_));
 sky130_fd_sc_hd__nand2_1 _17433_ (.A(_09603_),
    .B(_09533_),
    .Y(_13004_));
 sky130_fd_sc_hd__nand2_1 _17434_ (.A(_09602_),
    .B(_09548_),
    .Y(_13005_));
 sky130_fd_sc_hd__and3_1 _17435_ (.A(_13004_),
    .B(_09126_),
    .C(_13005_),
    .X(_13006_));
 sky130_fd_sc_hd__nand3_1 _17436_ (.A(_12960_),
    .B(_09052_),
    .C(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__nand2_1 _17437_ (.A(_12972_),
    .B(_09548_),
    .Y(_13008_));
 sky130_fd_sc_hd__o21ai_1 _17438_ (.A1(_13007_),
    .A2(_12971_),
    .B1(_13008_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand2_1 _17439_ (.A(_13005_),
    .B(_09016_),
    .Y(_13009_));
 sky130_fd_sc_hd__o21a_1 _17440_ (.A1(_09016_),
    .A2(_13005_),
    .B1(_09127_),
    .X(_13010_));
 sky130_fd_sc_hd__nand3_1 _17441_ (.A(_12960_),
    .B(_13009_),
    .C(_13010_),
    .Y(_13011_));
 sky130_fd_sc_hd__nand2_1 _17442_ (.A(_12972_),
    .B(net1959),
    .Y(_13012_));
 sky130_fd_sc_hd__o21ai_1 _17443_ (.A1(_13011_),
    .A2(_12971_),
    .B1(_13012_),
    .Y(_00160_));
 sky130_fd_sc_hd__inv_2 _17444_ (.A(net3829),
    .Y(_13013_));
 sky130_fd_sc_hd__nor2_2 _17445_ (.A(_12960_),
    .B(_12825_),
    .Y(_13014_));
 sky130_fd_sc_hd__nand2_4 _17446_ (.A(_08978_),
    .B(_09133_),
    .Y(_13015_));
 sky130_fd_sc_hd__nor2_1 _17447_ (.A(\res_v_active[0] ),
    .B(\res_v_active[1] ),
    .Y(_13016_));
 sky130_fd_sc_hd__inv_2 _17448_ (.A(\res_v_active[2] ),
    .Y(_13017_));
 sky130_fd_sc_hd__nand2_1 _17449_ (.A(_13016_),
    .B(_13017_),
    .Y(_13018_));
 sky130_fd_sc_hd__or2_1 _17450_ (.A(\res_v_active[3] ),
    .B(_13018_),
    .X(_13019_));
 sky130_fd_sc_hd__nor2_1 _17451_ (.A(\res_v_active[4] ),
    .B(_13019_),
    .Y(_13020_));
 sky130_fd_sc_hd__inv_2 _17452_ (.A(_13020_),
    .Y(_13021_));
 sky130_fd_sc_hd__or2_1 _17453_ (.A(\res_v_active[5] ),
    .B(_13021_),
    .X(_13022_));
 sky130_fd_sc_hd__nor2_1 _17454_ (.A(\res_v_active[6] ),
    .B(_13022_),
    .Y(_13023_));
 sky130_fd_sc_hd__or3b_1 _17455_ (.A(\res_v_counter[7] ),
    .B(_13023_),
    .C_N(\res_v_active[7] ),
    .X(_13024_));
 sky130_fd_sc_hd__inv_2 _17456_ (.A(net3451),
    .Y(_13025_));
 sky130_fd_sc_hd__inv_2 _17457_ (.A(_13023_),
    .Y(_13026_));
 sky130_fd_sc_hd__nand2_1 _17458_ (.A(_13022_),
    .B(\res_v_active[6] ),
    .Y(_13027_));
 sky130_fd_sc_hd__nand2_1 _17459_ (.A(_13026_),
    .B(_13027_),
    .Y(_13028_));
 sky130_fd_sc_hd__or2_1 _17460_ (.A(_13025_),
    .B(_13028_),
    .X(_13029_));
 sky130_fd_sc_hd__inv_2 _17461_ (.A(net3836),
    .Y(_13030_));
 sky130_fd_sc_hd__a21o_1 _17462_ (.A1(_13026_),
    .A2(\res_v_active[7] ),
    .B1(_13030_),
    .X(_13031_));
 sky130_fd_sc_hd__and3_1 _17463_ (.A(_13024_),
    .B(_13029_),
    .C(_13031_),
    .X(_13032_));
 sky130_fd_sc_hd__nand2_1 _17464_ (.A(_13019_),
    .B(\res_v_active[4] ),
    .Y(_13033_));
 sky130_fd_sc_hd__nand2_1 _17465_ (.A(_13021_),
    .B(_13033_),
    .Y(_13034_));
 sky130_fd_sc_hd__xor2_1 _17466_ (.A(\res_v_counter[4] ),
    .B(_13034_),
    .X(_13035_));
 sky130_fd_sc_hd__nand2_1 _17467_ (.A(_13018_),
    .B(\res_v_active[3] ),
    .Y(_13036_));
 sky130_fd_sc_hd__nand2_1 _17468_ (.A(_13019_),
    .B(_13036_),
    .Y(_13037_));
 sky130_fd_sc_hd__xnor2_1 _17469_ (.A(\res_v_counter[1] ),
    .B(\res_v_active[1] ),
    .Y(_13038_));
 sky130_fd_sc_hd__nand2_1 _17470_ (.A(_13013_),
    .B(\res_v_active[0] ),
    .Y(_13039_));
 sky130_fd_sc_hd__o21ai_1 _17471_ (.A1(\res_v_active[0] ),
    .A2(_13038_),
    .B1(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__o211ai_1 _17472_ (.A1(\res_v_counter[0] ),
    .A2(_13038_),
    .B1(_12323_),
    .C1(_13040_),
    .Y(_13041_));
 sky130_fd_sc_hd__or2_1 _17473_ (.A(_13017_),
    .B(_13016_),
    .X(_13042_));
 sky130_fd_sc_hd__nand2_1 _17474_ (.A(_13042_),
    .B(_13018_),
    .Y(_13043_));
 sky130_fd_sc_hd__nand2_1 _17475_ (.A(_13043_),
    .B(\res_v_counter[2] ),
    .Y(_13044_));
 sky130_fd_sc_hd__or2_1 _17476_ (.A(\res_v_counter[2] ),
    .B(_13043_),
    .X(_13045_));
 sky130_fd_sc_hd__a2bb2o_1 _17477_ (.A1_N(_12320_),
    .A2_N(_13037_),
    .B1(_13044_),
    .B2(_13045_),
    .X(_13046_));
 sky130_fd_sc_hd__a211o_1 _17478_ (.A1(_12320_),
    .A2(_13037_),
    .B1(_13041_),
    .C1(_13046_),
    .X(_13047_));
 sky130_fd_sc_hd__nor2_1 _17479_ (.A(_13035_),
    .B(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__nand2_1 _17480_ (.A(_13021_),
    .B(\res_v_active[5] ),
    .Y(_13049_));
 sky130_fd_sc_hd__nand2_1 _17481_ (.A(_13022_),
    .B(_13049_),
    .Y(_13050_));
 sky130_fd_sc_hd__inv_2 _17482_ (.A(net3777),
    .Y(_13051_));
 sky130_fd_sc_hd__nand2_1 _17483_ (.A(_13050_),
    .B(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__or2_1 _17484_ (.A(_13051_),
    .B(_13050_),
    .X(_13053_));
 sky130_fd_sc_hd__o211a_1 _17485_ (.A1(\res_v_active[7] ),
    .A2(_13026_),
    .B1(_13052_),
    .C1(_13053_),
    .X(_13054_));
 sky130_fd_sc_hd__nand2_1 _17486_ (.A(_13028_),
    .B(_13025_),
    .Y(_13055_));
 sky130_fd_sc_hd__and4_2 _17487_ (.A(_13032_),
    .B(_13048_),
    .C(_13054_),
    .D(_13055_),
    .X(_13056_));
 sky130_fd_sc_hd__nor2_1 _17488_ (.A(_13056_),
    .B(_13015_),
    .Y(_13057_));
 sky130_fd_sc_hd__or2_1 _17489_ (.A(net3829),
    .B(_13057_),
    .X(_13058_));
 sky130_fd_sc_hd__o2111ai_1 _17490_ (.A1(_13013_),
    .A2(_13015_),
    .B1(_09516_),
    .C1(_09114_),
    .D1(_13058_),
    .Y(_13059_));
 sky130_fd_sc_hd__o22ai_1 _17491_ (.A1(_13013_),
    .A2(_09497_),
    .B1(_13014_),
    .B2(_13059_),
    .Y(_00161_));
 sky130_fd_sc_hd__xor2_1 _17492_ (.A(_08829_),
    .B(_08830_),
    .X(_13060_));
 sky130_fd_sc_hd__xor2_1 _17493_ (.A(_09504_),
    .B(_13060_),
    .X(_13061_));
 sky130_fd_sc_hd__xor2_1 _17494_ (.A(\prescaler[3] ),
    .B(_08838_),
    .X(_13062_));
 sky130_fd_sc_hd__xor2_1 _17495_ (.A(_08836_),
    .B(_13062_),
    .X(_13063_));
 sky130_fd_sc_hd__or3_1 _17496_ (.A(_13061_),
    .B(_13063_),
    .C(_08846_),
    .X(_13064_));
 sky130_fd_sc_hd__and3_1 _17497_ (.A(_08830_),
    .B(_08829_),
    .C(_08831_),
    .X(_13065_));
 sky130_fd_sc_hd__clkbuf_2 _17498_ (.A(_13065_),
    .X(_13066_));
 sky130_fd_sc_hd__or2_1 _17499_ (.A(\prescaler_counter[8] ),
    .B(_13066_),
    .X(_13067_));
 sky130_fd_sc_hd__xor2_1 _17500_ (.A(\prescaler_counter[7] ),
    .B(_13066_),
    .X(_13068_));
 sky130_fd_sc_hd__xor2_1 _17501_ (.A(\prescaler_counter[6] ),
    .B(_13066_),
    .X(_13069_));
 sky130_fd_sc_hd__xor2_1 _17502_ (.A(\prescaler_counter[5] ),
    .B(_13066_),
    .X(_13070_));
 sky130_fd_sc_hd__xor2_1 _17503_ (.A(\prescaler_counter[4] ),
    .B(_13066_),
    .X(_13071_));
 sky130_fd_sc_hd__or4_1 _17504_ (.A(_13068_),
    .B(_13069_),
    .C(_13070_),
    .D(_13071_),
    .X(_13072_));
 sky130_fd_sc_hd__or4_1 _17505_ (.A(_09056_),
    .B(_13064_),
    .C(_13067_),
    .D(_13072_),
    .X(_13073_));
 sky130_fd_sc_hd__buf_2 _17506_ (.A(_13073_),
    .X(_13074_));
 sky130_fd_sc_hd__nand2_1 _17507_ (.A(net2003),
    .B(\res_v_counter[0] ),
    .Y(_13075_));
 sky130_fd_sc_hd__inv_2 _17508_ (.A(_13075_),
    .Y(_13076_));
 sky130_fd_sc_hd__nor2_1 _17509_ (.A(_12319_),
    .B(_13076_),
    .Y(_13077_));
 sky130_fd_sc_hd__a22o_1 _17510_ (.A1(net2003),
    .A2(_13015_),
    .B1(_13057_),
    .B2(_13077_),
    .X(_13078_));
 sky130_fd_sc_hd__nand2b_1 _17511_ (.A_N(_13074_),
    .B(_13078_),
    .Y(_13079_));
 sky130_fd_sc_hd__nand2_1 _17512_ (.A(_09498_),
    .B(net2003),
    .Y(_13080_));
 sky130_fd_sc_hd__o21ai_1 _17513_ (.A1(_13014_),
    .A2(_13079_),
    .B1(_13080_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _17514_ (.A(_12774_),
    .B(_12809_),
    .Y(_13081_));
 sky130_fd_sc_hd__nor3_1 _17515_ (.A(_13081_),
    .B(_12820_),
    .C(_12766_),
    .Y(_13082_));
 sky130_fd_sc_hd__nand2b_1 _17516_ (.A_N(_12823_),
    .B(_12814_),
    .Y(_13083_));
 sky130_fd_sc_hd__inv_2 _17517_ (.A(_13083_),
    .Y(_13084_));
 sky130_fd_sc_hd__nand3b_4 _17518_ (.A_N(_12960_),
    .B(_13082_),
    .C(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__xor2_1 _17519_ (.A(net3804),
    .B(_13075_),
    .X(_13086_));
 sky130_fd_sc_hd__or3_1 _17520_ (.A(_13056_),
    .B(_13086_),
    .C(_13015_),
    .X(_13087_));
 sky130_fd_sc_hd__nand2_1 _17521_ (.A(_13015_),
    .B(net3804),
    .Y(_13088_));
 sky130_fd_sc_hd__a21oi_1 _17522_ (.A1(_13087_),
    .A2(_13088_),
    .B1(_13074_),
    .Y(_02733_));
 sky130_fd_sc_hd__nand2_1 _17523_ (.A(_13085_),
    .B(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hd__o21ai_1 _17524_ (.A1(_12321_),
    .A2(_12682_),
    .B1(_02734_),
    .Y(_00163_));
 sky130_fd_sc_hd__and3_1 _17525_ (.A(_13076_),
    .B(net3749),
    .C(\res_v_counter[2] ),
    .X(_02735_));
 sky130_fd_sc_hd__o21ai_1 _17526_ (.A1(_12321_),
    .A2(_13075_),
    .B1(_12320_),
    .Y(_02736_));
 sky130_fd_sc_hd__or2b_1 _17527_ (.A(_02735_),
    .B_N(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__or3_1 _17528_ (.A(_13056_),
    .B(_02737_),
    .C(_13015_),
    .X(_02738_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_13015_),
    .B(net3749),
    .Y(_02739_));
 sky130_fd_sc_hd__a21oi_1 _17530_ (.A1(_02738_),
    .A2(_02739_),
    .B1(_13074_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_13085_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__o21ai_1 _17532_ (.A1(_12320_),
    .A2(_12682_),
    .B1(_02741_),
    .Y(_00164_));
 sky130_fd_sc_hd__or2_1 _17533_ (.A(net2497),
    .B(_02735_),
    .X(_02742_));
 sky130_fd_sc_hd__nand2_1 _17534_ (.A(_02735_),
    .B(net2497),
    .Y(_02743_));
 sky130_fd_sc_hd__and2_1 _17535_ (.A(_02742_),
    .B(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__a22o_1 _17536_ (.A1(net2497),
    .A2(_13015_),
    .B1(_13057_),
    .B2(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__nand2b_1 _17537_ (.A_N(_13074_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand2_1 _17538_ (.A(_09498_),
    .B(net2497),
    .Y(_02747_));
 sky130_fd_sc_hd__o21ai_1 _17539_ (.A1(_13014_),
    .A2(_02746_),
    .B1(_02747_),
    .Y(_00165_));
 sky130_fd_sc_hd__or2_1 _17540_ (.A(_13051_),
    .B(_02743_),
    .X(_02748_));
 sky130_fd_sc_hd__nand2_1 _17541_ (.A(_02743_),
    .B(_13051_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_1 _17542_ (.A(_02748_),
    .B(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__or3_1 _17543_ (.A(_13056_),
    .B(_02750_),
    .C(_13015_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_1 _17544_ (.A(_13015_),
    .B(net3777),
    .Y(_02752_));
 sky130_fd_sc_hd__a21oi_1 _17545_ (.A1(_02751_),
    .A2(_02752_),
    .B1(_13074_),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _17546_ (.A(_13085_),
    .B(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__o21ai_1 _17547_ (.A1(_13051_),
    .A2(_12682_),
    .B1(_02754_),
    .Y(_00166_));
 sky130_fd_sc_hd__or2_1 _17548_ (.A(_02748_),
    .B(_13015_),
    .X(_02755_));
 sky130_fd_sc_hd__or2_1 _17549_ (.A(_13025_),
    .B(_02748_),
    .X(_02756_));
 sky130_fd_sc_hd__or2b_1 _17550_ (.A(_13056_),
    .B_N(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__a31o_1 _17551_ (.A1(_08978_),
    .A2(_09133_),
    .A3(_02757_),
    .B1(_13074_),
    .X(_02758_));
 sky130_fd_sc_hd__a21o_1 _17552_ (.A1(_13025_),
    .A2(_02755_),
    .B1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__o22ai_1 _17553_ (.A1(_13025_),
    .A2(_09497_),
    .B1(_02759_),
    .B2(_13014_),
    .Y(_00167_));
 sky130_fd_sc_hd__or2_1 _17554_ (.A(_02756_),
    .B(_13015_),
    .X(_02760_));
 sky130_fd_sc_hd__or2_1 _17555_ (.A(_13030_),
    .B(_02756_),
    .X(_02761_));
 sky130_fd_sc_hd__or2b_1 _17556_ (.A(_13056_),
    .B_N(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__a31o_1 _17557_ (.A1(_08978_),
    .A2(_09133_),
    .A3(_02762_),
    .B1(_13074_),
    .X(_02763_));
 sky130_fd_sc_hd__a21o_1 _17558_ (.A1(_13030_),
    .A2(_02760_),
    .B1(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__o22ai_1 _17559_ (.A1(_13030_),
    .A2(_09497_),
    .B1(_02764_),
    .B2(_13014_),
    .Y(_00168_));
 sky130_fd_sc_hd__inv_2 _17560_ (.A(net2028),
    .Y(_02765_));
 sky130_fd_sc_hd__or2_1 _17561_ (.A(_02761_),
    .B(_13015_),
    .X(_02766_));
 sky130_fd_sc_hd__or2_1 _17562_ (.A(_02765_),
    .B(_02761_),
    .X(_02767_));
 sky130_fd_sc_hd__or2b_1 _17563_ (.A(_13056_),
    .B_N(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__a31o_1 _17564_ (.A1(_08978_),
    .A2(_09133_),
    .A3(_02768_),
    .B1(_13074_),
    .X(_02769_));
 sky130_fd_sc_hd__a21o_1 _17565_ (.A1(_02765_),
    .A2(_02766_),
    .B1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__o22ai_1 _17566_ (.A1(_02765_),
    .A2(_09497_),
    .B1(_02770_),
    .B2(_13014_),
    .Y(_00169_));
 sky130_fd_sc_hd__nor2_1 _17567_ (.A(_08992_),
    .B(_02767_),
    .Y(_02771_));
 sky130_fd_sc_hd__xnor2_1 _17568_ (.A(net2057),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__or2_1 _17569_ (.A(_02772_),
    .B(_09119_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_1 _17570_ (.A(_09119_),
    .B(net2057),
    .Y(_02774_));
 sky130_fd_sc_hd__a21oi_1 _17571_ (.A1(_02773_),
    .A2(_02774_),
    .B1(_13074_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_1 _17572_ (.A(_13085_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__nand2_1 _17573_ (.A(_09498_),
    .B(net2057),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _17574_ (.A(_02776_),
    .B(_02777_),
    .Y(_00170_));
 sky130_fd_sc_hd__nor2_1 _17575_ (.A(net2014),
    .B(_12968_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand2_1 _17576_ (.A(_12960_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__nand2_2 _17577_ (.A(_12966_),
    .B(_09497_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_1 _17578_ (.A(_02780_),
    .B(net2014),
    .Y(_02781_));
 sky130_fd_sc_hd__o21ai_1 _17579_ (.A1(_02779_),
    .A2(_02780_),
    .B1(net2015),
    .Y(_00171_));
 sky130_fd_sc_hd__nand2_1 _17580_ (.A(\pixel_double_counter[0] ),
    .B(net1999),
    .Y(_02782_));
 sky130_fd_sc_hd__or2_1 _17581_ (.A(\pixel_double_counter[0] ),
    .B(net1999),
    .X(_02783_));
 sky130_fd_sc_hd__and3_1 _17582_ (.A(_12967_),
    .B(_02782_),
    .C(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__nand2_1 _17583_ (.A(_12960_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__nand2_1 _17584_ (.A(_02780_),
    .B(net1999),
    .Y(_02786_));
 sky130_fd_sc_hd__o21ai_1 _17585_ (.A1(_02785_),
    .A2(_02780_),
    .B1(net2000),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _17586_ (.A(_02782_),
    .B(_08865_),
    .Y(_02787_));
 sky130_fd_sc_hd__or2_1 _17587_ (.A(_08865_),
    .B(_02782_),
    .X(_02788_));
 sky130_fd_sc_hd__and3_1 _17588_ (.A(_12967_),
    .B(_02787_),
    .C(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__nand2_1 _17589_ (.A(_12960_),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__nand2_1 _17590_ (.A(_02780_),
    .B(net1940),
    .Y(_02791_));
 sky130_fd_sc_hd__o21ai_1 _17591_ (.A1(_02790_),
    .A2(_02780_),
    .B1(net1941),
    .Y(_00173_));
 sky130_fd_sc_hd__a21oi_1 _17592_ (.A1(_02788_),
    .A2(_08861_),
    .B1(_12851_),
    .Y(_02792_));
 sky130_fd_sc_hd__o211a_1 _17593_ (.A1(_08861_),
    .A2(_02788_),
    .B1(_02792_),
    .C1(_08870_),
    .X(_02793_));
 sky130_fd_sc_hd__nand2_1 _17594_ (.A(_12960_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__nand2_1 _17595_ (.A(_02780_),
    .B(net1862),
    .Y(_02795_));
 sky130_fd_sc_hd__o21ai_1 _17596_ (.A1(_02794_),
    .A2(_02780_),
    .B1(net1863),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _17597_ (.A(_08992_),
    .B(_09126_),
    .Y(_02796_));
 sky130_fd_sc_hd__or2_1 _17598_ (.A(net2110),
    .B(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__nand2_1 _17599_ (.A(_08980_),
    .B(_09052_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_2 _17600_ (.A(_02798_),
    .B(_09058_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand2_1 _17601_ (.A(_02799_),
    .B(net2110),
    .Y(_02800_));
 sky130_fd_sc_hd__o21ai_1 _17602_ (.A1(_02797_),
    .A2(_02799_),
    .B1(net2111),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _17603_ (.A(_08981_),
    .B(net2110),
    .Y(_02801_));
 sky130_fd_sc_hd__or2_1 _17604_ (.A(_02796_),
    .B(_02799_),
    .X(_02802_));
 sky130_fd_sc_hd__a31o_1 _17605_ (.A1(_02798_),
    .A2(_09058_),
    .A3(_02797_),
    .B1(_08981_),
    .X(_02803_));
 sky130_fd_sc_hd__o21ai_1 _17606_ (.A1(_02801_),
    .A2(_02802_),
    .B1(_02803_),
    .Y(_00176_));
 sky130_fd_sc_hd__or3b_1 _17607_ (.A(_08981_),
    .B(_08986_),
    .C_N(\line_double_counter[0] ),
    .X(_02804_));
 sky130_fd_sc_hd__a21o_1 _17608_ (.A1(\line_double_counter[0] ),
    .A2(\line_double_counter[1] ),
    .B1(net1992),
    .X(_02805_));
 sky130_fd_sc_hd__nand2_1 _17609_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__o2bb2ai_1 _17610_ (.A1_N(net1992),
    .A2_N(_02799_),
    .B1(_02806_),
    .B2(_02802_),
    .Y(_00177_));
 sky130_fd_sc_hd__xor2_1 _17611_ (.A(net2005),
    .B(_02804_),
    .X(_02807_));
 sky130_fd_sc_hd__o2bb2ai_1 _17612_ (.A1_N(net2005),
    .A2_N(_02799_),
    .B1(_02807_),
    .B2(_02802_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _17613_ (.A(_09126_),
    .B(_12183_),
    .Y(_02808_));
 sky130_fd_sc_hd__clkinv_4 _17614_ (.A(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__buf_8 _17615_ (.A(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__nor2_1 _17616_ (.A(\line_cache_idx[3] ),
    .B(\line_cache_idx[2] ),
    .Y(_02811_));
 sky130_fd_sc_hd__clkinv_4 _17617_ (.A(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__nor2_2 _17618_ (.A(\line_cache_idx[4] ),
    .B(\line_cache_idx[5] ),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_2 _17619_ (.A(_12174_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__nor2_1 _17620_ (.A(_02812_),
    .B(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__inv_2 _17621_ (.A(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__nor2_2 _17622_ (.A(_12177_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__clkbuf_16 _17623_ (.A(_12190_),
    .X(_02818_));
 sky130_fd_sc_hd__o21ai_4 _17624_ (.A1(_12290_),
    .A2(_02817_),
    .B1(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__mux2_1 _17625_ (.A0(_02810_),
    .A1(net2260),
    .S(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _17626_ (.A(_02820_),
    .X(_00179_));
 sky130_fd_sc_hd__nand2_1 _17627_ (.A(_09126_),
    .B(_12196_),
    .Y(_02821_));
 sky130_fd_sc_hd__clkinv_4 _17628_ (.A(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__buf_8 _17629_ (.A(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__mux2_1 _17630_ (.A0(_02823_),
    .A1(net2020),
    .S(_02819_),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_1 _17631_ (.A(_02824_),
    .X(_00180_));
 sky130_fd_sc_hd__nand2_1 _17632_ (.A(_12180_),
    .B(_12204_),
    .Y(_02825_));
 sky130_fd_sc_hd__clkinv_4 _17633_ (.A(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__buf_8 _17634_ (.A(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _17635_ (.A0(_02827_),
    .A1(net2362),
    .S(_02819_),
    .X(_02828_));
 sky130_fd_sc_hd__clkbuf_1 _17636_ (.A(_02828_),
    .X(_00181_));
 sky130_fd_sc_hd__nand2_1 _17637_ (.A(_12180_),
    .B(_12212_),
    .Y(_02829_));
 sky130_fd_sc_hd__clkinv_4 _17638_ (.A(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__buf_8 _17639_ (.A(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _17640_ (.A0(_02831_),
    .A1(net2050),
    .S(_02819_),
    .X(_02832_));
 sky130_fd_sc_hd__clkbuf_1 _17641_ (.A(_02832_),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_1 _17642_ (.A(_12180_),
    .B(_12220_),
    .Y(_02833_));
 sky130_fd_sc_hd__clkinv_4 _17643_ (.A(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__clkbuf_16 _17644_ (.A(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _17645_ (.A0(_02835_),
    .A1(net3434),
    .S(_02819_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _17646_ (.A(_02836_),
    .X(_00183_));
 sky130_fd_sc_hd__nand2_1 _17647_ (.A(_12180_),
    .B(_12228_),
    .Y(_02837_));
 sky130_fd_sc_hd__inv_4 _17648_ (.A(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__buf_8 _17649_ (.A(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__mux2_1 _17650_ (.A0(_02839_),
    .A1(net2912),
    .S(_02819_),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _17651_ (.A(_02840_),
    .X(_00184_));
 sky130_fd_sc_hd__nand2_1 _17652_ (.A(_12180_),
    .B(_12236_),
    .Y(_02841_));
 sky130_fd_sc_hd__clkinv_4 _17653_ (.A(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__buf_8 _17654_ (.A(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _17655_ (.A0(_02843_),
    .A1(net2348),
    .S(_02819_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _17656_ (.A(_02844_),
    .X(_00185_));
 sky130_fd_sc_hd__nand2_1 _17657_ (.A(_12180_),
    .B(_12244_),
    .Y(_02845_));
 sky130_fd_sc_hd__clkinv_4 _17658_ (.A(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__buf_8 _17659_ (.A(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(_02847_),
    .A1(net2887),
    .S(_02819_),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _17661_ (.A(_02848_),
    .X(_00186_));
 sky130_fd_sc_hd__buf_4 _17662_ (.A(_02819_),
    .X(_02849_));
 sky130_fd_sc_hd__buf_12 _17663_ (.A(net81),
    .X(_02850_));
 sky130_fd_sc_hd__inv_2 _17664_ (.A(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__buf_8 _17665_ (.A(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__buf_4 _17666_ (.A(_02817_),
    .X(_02853_));
 sky130_fd_sc_hd__buf_8 _17667_ (.A(_12183_),
    .X(_02854_));
 sky130_fd_sc_hd__buf_4 _17668_ (.A(_02817_),
    .X(_02855_));
 sky130_fd_sc_hd__nor2_1 _17669_ (.A(_02854_),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__a211o_1 _17670_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__buf_4 _17671_ (.A(_02819_),
    .X(_02858_));
 sky130_fd_sc_hd__nand2_1 _17672_ (.A(_02858_),
    .B(net430),
    .Y(_02859_));
 sky130_fd_sc_hd__o21ai_1 _17673_ (.A1(_02849_),
    .A2(_02857_),
    .B1(net431),
    .Y(_00187_));
 sky130_fd_sc_hd__buf_12 _17674_ (.A(net82),
    .X(_02860_));
 sky130_fd_sc_hd__inv_2 _17675_ (.A(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__clkbuf_16 _17676_ (.A(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_16 _17677_ (.A(_12196_),
    .X(_02863_));
 sky130_fd_sc_hd__nor2_1 _17678_ (.A(_02863_),
    .B(_02855_),
    .Y(_02864_));
 sky130_fd_sc_hd__a211o_1 _17679_ (.A1(_02862_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _17680_ (.A(_02858_),
    .B(net424),
    .Y(_02866_));
 sky130_fd_sc_hd__o21ai_1 _17681_ (.A1(_02849_),
    .A2(_02865_),
    .B1(net425),
    .Y(_00188_));
 sky130_fd_sc_hd__buf_12 _17682_ (.A(net51),
    .X(_02867_));
 sky130_fd_sc_hd__clkinv_4 _17683_ (.A(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__clkbuf_16 _17684_ (.A(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__buf_12 _17685_ (.A(_12204_),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_1 _17686_ (.A(_02870_),
    .B(_02855_),
    .Y(_02871_));
 sky130_fd_sc_hd__a211o_1 _17687_ (.A1(_02869_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__nand2_1 _17688_ (.A(_02858_),
    .B(net792),
    .Y(_02873_));
 sky130_fd_sc_hd__o21ai_1 _17689_ (.A1(_02849_),
    .A2(_02872_),
    .B1(net793),
    .Y(_00189_));
 sky130_fd_sc_hd__buf_12 _17690_ (.A(net52),
    .X(_02874_));
 sky130_fd_sc_hd__inv_2 _17691_ (.A(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__clkbuf_16 _17692_ (.A(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_16 _17693_ (.A(_12212_),
    .X(_02877_));
 sky130_fd_sc_hd__nor2_1 _17694_ (.A(_02877_),
    .B(_02855_),
    .Y(_02878_));
 sky130_fd_sc_hd__a211o_1 _17695_ (.A1(_02876_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__nand2_1 _17696_ (.A(_02858_),
    .B(net436),
    .Y(_02880_));
 sky130_fd_sc_hd__o21ai_1 _17697_ (.A1(_02849_),
    .A2(_02879_),
    .B1(net437),
    .Y(_00190_));
 sky130_fd_sc_hd__buf_12 _17698_ (.A(net53),
    .X(_02881_));
 sky130_fd_sc_hd__clkinv_4 _17699_ (.A(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__buf_12 _17700_ (.A(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_16 _17701_ (.A(_12220_),
    .X(_02884_));
 sky130_fd_sc_hd__nor2_1 _17702_ (.A(_02884_),
    .B(_02855_),
    .Y(_02885_));
 sky130_fd_sc_hd__a211o_1 _17703_ (.A1(_02883_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__nand2_1 _17704_ (.A(_02858_),
    .B(net534),
    .Y(_02887_));
 sky130_fd_sc_hd__o21ai_1 _17705_ (.A1(_02849_),
    .A2(_02886_),
    .B1(net535),
    .Y(_00191_));
 sky130_fd_sc_hd__buf_12 _17706_ (.A(net54),
    .X(_02888_));
 sky130_fd_sc_hd__clkinv_4 _17707_ (.A(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__buf_8 _17708_ (.A(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__clkbuf_16 _17709_ (.A(_12228_),
    .X(_02891_));
 sky130_fd_sc_hd__nor2_1 _17710_ (.A(_02891_),
    .B(_02855_),
    .Y(_02892_));
 sky130_fd_sc_hd__a211o_1 _17711_ (.A1(_02890_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_1 _17712_ (.A(_02858_),
    .B(net778),
    .Y(_02894_));
 sky130_fd_sc_hd__o21ai_1 _17713_ (.A1(_02849_),
    .A2(_02893_),
    .B1(net779),
    .Y(_00192_));
 sky130_fd_sc_hd__buf_12 _17714_ (.A(net55),
    .X(_02895_));
 sky130_fd_sc_hd__clkinv_4 _17715_ (.A(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__buf_12 _17716_ (.A(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_16 _17717_ (.A(_12236_),
    .X(_02898_));
 sky130_fd_sc_hd__nor2_1 _17718_ (.A(_02898_),
    .B(_02855_),
    .Y(_02899_));
 sky130_fd_sc_hd__a211o_1 _17719_ (.A1(_02897_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__nand2_1 _17720_ (.A(_02858_),
    .B(net466),
    .Y(_02901_));
 sky130_fd_sc_hd__o21ai_1 _17721_ (.A1(_02849_),
    .A2(_02900_),
    .B1(net467),
    .Y(_00193_));
 sky130_fd_sc_hd__clkbuf_16 _17722_ (.A(net56),
    .X(_02902_));
 sky130_fd_sc_hd__clkinv_4 _17723_ (.A(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__clkbuf_16 _17724_ (.A(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__clkbuf_16 _17725_ (.A(_12244_),
    .X(_02905_));
 sky130_fd_sc_hd__nor2_1 _17726_ (.A(_02905_),
    .B(_02855_),
    .Y(_02906_));
 sky130_fd_sc_hd__a211o_1 _17727_ (.A1(_02904_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__nand2_1 _17728_ (.A(_02858_),
    .B(net406),
    .Y(_02908_));
 sky130_fd_sc_hd__o21ai_1 _17729_ (.A1(_02849_),
    .A2(_02907_),
    .B1(net407),
    .Y(_00194_));
 sky130_fd_sc_hd__buf_4 _17730_ (.A(_02819_),
    .X(_02909_));
 sky130_fd_sc_hd__buf_12 _17731_ (.A(net57),
    .X(_02910_));
 sky130_fd_sc_hd__inv_2 _17732_ (.A(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__buf_8 _17733_ (.A(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__a211o_1 _17734_ (.A1(_02912_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02856_),
    .X(_02913_));
 sky130_fd_sc_hd__nand2_1 _17735_ (.A(_02858_),
    .B(net530),
    .Y(_02914_));
 sky130_fd_sc_hd__o21ai_1 _17736_ (.A1(_02909_),
    .A2(_02913_),
    .B1(net531),
    .Y(_00195_));
 sky130_fd_sc_hd__buf_12 _17737_ (.A(net58),
    .X(_02915_));
 sky130_fd_sc_hd__clkinv_4 _17738_ (.A(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__clkbuf_16 _17739_ (.A(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__a211o_1 _17740_ (.A1(_02917_),
    .A2(_02853_),
    .B1(_09130_),
    .C1(_02864_),
    .X(_02918_));
 sky130_fd_sc_hd__nand2_1 _17741_ (.A(_02858_),
    .B(net904),
    .Y(_02919_));
 sky130_fd_sc_hd__o21ai_1 _17742_ (.A1(_02909_),
    .A2(_02918_),
    .B1(net905),
    .Y(_00196_));
 sky130_fd_sc_hd__buf_12 _17743_ (.A(net59),
    .X(_02920_));
 sky130_fd_sc_hd__clkinv_4 _17744_ (.A(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__clkbuf_16 _17745_ (.A(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__buf_4 _17746_ (.A(_09129_),
    .X(_02923_));
 sky130_fd_sc_hd__a211o_1 _17747_ (.A1(_02922_),
    .A2(_02853_),
    .B1(_02923_),
    .C1(_02871_),
    .X(_02924_));
 sky130_fd_sc_hd__nand2_1 _17748_ (.A(_02858_),
    .B(net470),
    .Y(_02925_));
 sky130_fd_sc_hd__o21ai_1 _17749_ (.A1(_02909_),
    .A2(_02924_),
    .B1(net471),
    .Y(_00197_));
 sky130_fd_sc_hd__buf_12 _17750_ (.A(net60),
    .X(_02926_));
 sky130_fd_sc_hd__clkinv_4 _17751_ (.A(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__clkbuf_16 _17752_ (.A(_02927_),
    .X(_02928_));
 sky130_fd_sc_hd__a211o_1 _17753_ (.A1(_02928_),
    .A2(_02853_),
    .B1(_02923_),
    .C1(_02878_),
    .X(_02929_));
 sky130_fd_sc_hd__nand2_1 _17754_ (.A(_02858_),
    .B(net452),
    .Y(_02930_));
 sky130_fd_sc_hd__o21ai_1 _17755_ (.A1(_02909_),
    .A2(_02929_),
    .B1(net453),
    .Y(_00198_));
 sky130_fd_sc_hd__buf_12 _17756_ (.A(net62),
    .X(_02931_));
 sky130_fd_sc_hd__clkinv_4 _17757_ (.A(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__clkbuf_16 _17758_ (.A(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a211o_1 _17759_ (.A1(_02933_),
    .A2(_02853_),
    .B1(_02923_),
    .C1(_02885_),
    .X(_02934_));
 sky130_fd_sc_hd__nand2_1 _17760_ (.A(_02858_),
    .B(net414),
    .Y(_02935_));
 sky130_fd_sc_hd__o21ai_1 _17761_ (.A1(_02909_),
    .A2(_02934_),
    .B1(net415),
    .Y(_00199_));
 sky130_fd_sc_hd__buf_12 _17762_ (.A(net63),
    .X(_02936_));
 sky130_fd_sc_hd__clkinv_4 _17763_ (.A(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__buf_8 _17764_ (.A(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__a211o_1 _17765_ (.A1(_02938_),
    .A2(_02853_),
    .B1(_02923_),
    .C1(_02892_),
    .X(_02939_));
 sky130_fd_sc_hd__nand2_1 _17766_ (.A(_02858_),
    .B(net440),
    .Y(_02940_));
 sky130_fd_sc_hd__o21ai_1 _17767_ (.A1(_02909_),
    .A2(_02939_),
    .B1(net441),
    .Y(_00200_));
 sky130_fd_sc_hd__buf_12 _17768_ (.A(net64),
    .X(_02941_));
 sky130_fd_sc_hd__clkinv_4 _17769_ (.A(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__buf_12 _17770_ (.A(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__a211o_1 _17771_ (.A1(_02943_),
    .A2(_02853_),
    .B1(_02923_),
    .C1(_02899_),
    .X(_02944_));
 sky130_fd_sc_hd__nand2_1 _17772_ (.A(_02858_),
    .B(net398),
    .Y(_02945_));
 sky130_fd_sc_hd__o21ai_1 _17773_ (.A1(_02909_),
    .A2(_02944_),
    .B1(net399),
    .Y(_00201_));
 sky130_fd_sc_hd__clkbuf_16 _17774_ (.A(net65),
    .X(_02946_));
 sky130_fd_sc_hd__clkinv_4 _17775_ (.A(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__clkbuf_16 _17776_ (.A(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__a211o_1 _17777_ (.A1(_02948_),
    .A2(_02853_),
    .B1(_02923_),
    .C1(_02906_),
    .X(_02949_));
 sky130_fd_sc_hd__nand2_1 _17778_ (.A(_02858_),
    .B(net608),
    .Y(_02950_));
 sky130_fd_sc_hd__o21ai_1 _17779_ (.A1(_02909_),
    .A2(_02949_),
    .B1(net609),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _17780_ (.A(_12169_),
    .Y(_02951_));
 sky130_fd_sc_hd__buf_8 _17781_ (.A(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__a211o_1 _17782_ (.A1(_02952_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02856_),
    .X(_02953_));
 sky130_fd_sc_hd__nand2_1 _17783_ (.A(_02849_),
    .B(net1352),
    .Y(_02954_));
 sky130_fd_sc_hd__o21ai_1 _17784_ (.A1(_02909_),
    .A2(_02953_),
    .B1(net1353),
    .Y(_00203_));
 sky130_fd_sc_hd__clkinv_4 _17785_ (.A(_12194_),
    .Y(_02955_));
 sky130_fd_sc_hd__clkbuf_16 _17786_ (.A(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__a211o_1 _17787_ (.A1(_02956_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02864_),
    .X(_02957_));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(_02849_),
    .B(net1840),
    .Y(_02958_));
 sky130_fd_sc_hd__o21ai_1 _17789_ (.A1(_02909_),
    .A2(_02957_),
    .B1(net1841),
    .Y(_00204_));
 sky130_fd_sc_hd__clkinv_4 _17790_ (.A(_12202_),
    .Y(_02959_));
 sky130_fd_sc_hd__clkbuf_16 _17791_ (.A(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__a211o_1 _17792_ (.A1(_02960_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02871_),
    .X(_02961_));
 sky130_fd_sc_hd__nand2_1 _17793_ (.A(_02849_),
    .B(net1962),
    .Y(_02962_));
 sky130_fd_sc_hd__o21ai_1 _17794_ (.A1(_02909_),
    .A2(_02961_),
    .B1(_02962_),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _17795_ (.A(_12210_),
    .Y(_02963_));
 sky130_fd_sc_hd__clkbuf_16 _17796_ (.A(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__a211o_1 _17797_ (.A1(_02964_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02878_),
    .X(_02965_));
 sky130_fd_sc_hd__nand2_1 _17798_ (.A(_02849_),
    .B(net1927),
    .Y(_02966_));
 sky130_fd_sc_hd__o21ai_1 _17799_ (.A1(_02909_),
    .A2(_02965_),
    .B1(net1928),
    .Y(_00206_));
 sky130_fd_sc_hd__clkinv_4 _17800_ (.A(_12218_),
    .Y(_02967_));
 sky130_fd_sc_hd__buf_12 _17801_ (.A(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__a211o_1 _17802_ (.A1(_02968_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02885_),
    .X(_02969_));
 sky130_fd_sc_hd__nand2_1 _17803_ (.A(_02849_),
    .B(net1950),
    .Y(_02970_));
 sky130_fd_sc_hd__o21ai_1 _17804_ (.A1(_02909_),
    .A2(_02969_),
    .B1(_02970_),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _17805_ (.A(_12226_),
    .Y(_02971_));
 sky130_fd_sc_hd__buf_8 _17806_ (.A(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__a211o_1 _17807_ (.A1(_02972_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02892_),
    .X(_02973_));
 sky130_fd_sc_hd__nand2_1 _17808_ (.A(_02849_),
    .B(net1881),
    .Y(_02974_));
 sky130_fd_sc_hd__o21ai_1 _17809_ (.A1(_02909_),
    .A2(_02973_),
    .B1(net1882),
    .Y(_00208_));
 sky130_fd_sc_hd__inv_2 _17810_ (.A(_12234_),
    .Y(_02975_));
 sky130_fd_sc_hd__buf_12 _17811_ (.A(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__a211o_1 _17812_ (.A1(_02976_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02899_),
    .X(_02977_));
 sky130_fd_sc_hd__nand2_1 _17813_ (.A(_02849_),
    .B(net1202),
    .Y(_02978_));
 sky130_fd_sc_hd__o21ai_1 _17814_ (.A1(_02909_),
    .A2(_02977_),
    .B1(net1203),
    .Y(_00209_));
 sky130_fd_sc_hd__clkinv_4 _17815_ (.A(_12242_),
    .Y(_02979_));
 sky130_fd_sc_hd__clkbuf_16 _17816_ (.A(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__a211o_1 _17817_ (.A1(_02980_),
    .A2(_02855_),
    .B1(_02923_),
    .C1(_02906_),
    .X(_02981_));
 sky130_fd_sc_hd__nand2_1 _17818_ (.A(_02849_),
    .B(net1072),
    .Y(_02982_));
 sky130_fd_sc_hd__o21ai_1 _17819_ (.A1(_02909_),
    .A2(_02981_),
    .B1(net1073),
    .Y(_00210_));
 sky130_fd_sc_hd__nor2_1 _17820_ (.A(_12293_),
    .B(_02814_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_1 _17821_ (.A(_02983_),
    .B(_12313_),
    .Y(_02984_));
 sky130_fd_sc_hd__inv_2 _17822_ (.A(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__o21ai_4 _17823_ (.A1(_12290_),
    .A2(_02985_),
    .B1(_02818_),
    .Y(_02986_));
 sky130_fd_sc_hd__mux2_1 _17824_ (.A0(_02810_),
    .A1(net2731),
    .S(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__clkbuf_1 _17825_ (.A(_02987_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _17826_ (.A0(_02823_),
    .A1(net2225),
    .S(_02986_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_1 _17827_ (.A(_02988_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _17828_ (.A0(_02827_),
    .A1(net2250),
    .S(_02986_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _17829_ (.A(_02989_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _17830_ (.A0(_02831_),
    .A1(net2192),
    .S(_02986_),
    .X(_02990_));
 sky130_fd_sc_hd__clkbuf_1 _17831_ (.A(_02990_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _17832_ (.A0(_02835_),
    .A1(net3073),
    .S(_02986_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _17833_ (.A(_02991_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _17834_ (.A0(_02839_),
    .A1(net2772),
    .S(_02986_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _17835_ (.A(_02992_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _17836_ (.A0(_02843_),
    .A1(net2336),
    .S(_02986_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _17837_ (.A(_02993_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _17838_ (.A0(_02847_),
    .A1(net2205),
    .S(_02986_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _17839_ (.A(_02994_),
    .X(_00218_));
 sky130_fd_sc_hd__buf_4 _17840_ (.A(_02986_),
    .X(_02995_));
 sky130_fd_sc_hd__buf_4 _17841_ (.A(_02985_),
    .X(_02996_));
 sky130_fd_sc_hd__buf_4 _17842_ (.A(_02985_),
    .X(_02997_));
 sky130_fd_sc_hd__nor2_1 _17843_ (.A(_02854_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__a211o_1 _17844_ (.A1(_02852_),
    .A2(_02996_),
    .B1(_02923_),
    .C1(_02998_),
    .X(_02999_));
 sky130_fd_sc_hd__buf_4 _17845_ (.A(_02986_),
    .X(_03000_));
 sky130_fd_sc_hd__nand2_1 _17846_ (.A(_03000_),
    .B(net956),
    .Y(_03001_));
 sky130_fd_sc_hd__o21ai_1 _17847_ (.A1(_02995_),
    .A2(_02999_),
    .B1(net957),
    .Y(_00219_));
 sky130_fd_sc_hd__nor2_1 _17848_ (.A(_02863_),
    .B(_02997_),
    .Y(_03002_));
 sky130_fd_sc_hd__a211o_1 _17849_ (.A1(_02862_),
    .A2(_02996_),
    .B1(_02923_),
    .C1(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__nand2_1 _17850_ (.A(_03000_),
    .B(net1254),
    .Y(_03004_));
 sky130_fd_sc_hd__o21ai_1 _17851_ (.A1(_02995_),
    .A2(_03003_),
    .B1(net1255),
    .Y(_00220_));
 sky130_fd_sc_hd__buf_4 _17852_ (.A(_09129_),
    .X(_03005_));
 sky130_fd_sc_hd__nor2_1 _17853_ (.A(_02870_),
    .B(_02997_),
    .Y(_03006_));
 sky130_fd_sc_hd__a211o_1 _17854_ (.A1(_02869_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__nand2_1 _17855_ (.A(_03000_),
    .B(net1586),
    .Y(_03008_));
 sky130_fd_sc_hd__o21ai_1 _17856_ (.A1(_02995_),
    .A2(_03007_),
    .B1(net1587),
    .Y(_00221_));
 sky130_fd_sc_hd__nor2_1 _17857_ (.A(_02877_),
    .B(_02997_),
    .Y(_03009_));
 sky130_fd_sc_hd__a211o_1 _17858_ (.A1(_02876_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__nand2_1 _17859_ (.A(_03000_),
    .B(net1186),
    .Y(_03011_));
 sky130_fd_sc_hd__o21ai_1 _17860_ (.A1(_02995_),
    .A2(_03010_),
    .B1(net1187),
    .Y(_00222_));
 sky130_fd_sc_hd__nor2_1 _17861_ (.A(_02884_),
    .B(_02997_),
    .Y(_03012_));
 sky130_fd_sc_hd__a211o_1 _17862_ (.A1(_02883_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__nand2_1 _17863_ (.A(_03000_),
    .B(net1694),
    .Y(_03014_));
 sky130_fd_sc_hd__o21ai_1 _17864_ (.A1(_02995_),
    .A2(_03013_),
    .B1(net1695),
    .Y(_00223_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(_02891_),
    .B(_02997_),
    .Y(_03015_));
 sky130_fd_sc_hd__a211o_1 _17866_ (.A1(_02890_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__nand2_1 _17867_ (.A(_03000_),
    .B(net814),
    .Y(_03017_));
 sky130_fd_sc_hd__o21ai_1 _17868_ (.A1(_02995_),
    .A2(_03016_),
    .B1(net815),
    .Y(_00224_));
 sky130_fd_sc_hd__nor2_1 _17869_ (.A(_02898_),
    .B(_02997_),
    .Y(_03018_));
 sky130_fd_sc_hd__a211o_1 _17870_ (.A1(_02897_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__nand2_1 _17871_ (.A(_03000_),
    .B(net948),
    .Y(_03020_));
 sky130_fd_sc_hd__o21ai_1 _17872_ (.A1(_02995_),
    .A2(_03019_),
    .B1(net949),
    .Y(_00225_));
 sky130_fd_sc_hd__nor2_1 _17873_ (.A(_02905_),
    .B(_02997_),
    .Y(_03021_));
 sky130_fd_sc_hd__a211o_1 _17874_ (.A1(_02904_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__nand2_1 _17875_ (.A(_03000_),
    .B(net1020),
    .Y(_03023_));
 sky130_fd_sc_hd__o21ai_1 _17876_ (.A1(_02995_),
    .A2(_03022_),
    .B1(net1021),
    .Y(_00226_));
 sky130_fd_sc_hd__buf_4 _17877_ (.A(_02986_),
    .X(_03024_));
 sky130_fd_sc_hd__a211o_1 _17878_ (.A1(_02912_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_02998_),
    .X(_03025_));
 sky130_fd_sc_hd__nand2_1 _17879_ (.A(_03000_),
    .B(net1828),
    .Y(_03026_));
 sky130_fd_sc_hd__o21ai_1 _17880_ (.A1(_03024_),
    .A2(_03025_),
    .B1(net1829),
    .Y(_00227_));
 sky130_fd_sc_hd__a211o_1 _17881_ (.A1(_02917_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03002_),
    .X(_03027_));
 sky130_fd_sc_hd__nand2_1 _17882_ (.A(_03000_),
    .B(net1328),
    .Y(_03028_));
 sky130_fd_sc_hd__o21ai_1 _17883_ (.A1(_03024_),
    .A2(_03027_),
    .B1(net1329),
    .Y(_00228_));
 sky130_fd_sc_hd__a211o_1 _17884_ (.A1(_02922_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03006_),
    .X(_03029_));
 sky130_fd_sc_hd__nand2_1 _17885_ (.A(_03000_),
    .B(net1802),
    .Y(_03030_));
 sky130_fd_sc_hd__o21ai_1 _17886_ (.A1(_03024_),
    .A2(_03029_),
    .B1(net1803),
    .Y(_00229_));
 sky130_fd_sc_hd__a211o_1 _17887_ (.A1(_02928_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03009_),
    .X(_03031_));
 sky130_fd_sc_hd__nand2_1 _17888_ (.A(_03000_),
    .B(net1664),
    .Y(_03032_));
 sky130_fd_sc_hd__o21ai_1 _17889_ (.A1(_03024_),
    .A2(_03031_),
    .B1(net1665),
    .Y(_00230_));
 sky130_fd_sc_hd__a211o_1 _17890_ (.A1(_02933_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03012_),
    .X(_03033_));
 sky130_fd_sc_hd__nand2_1 _17891_ (.A(_03000_),
    .B(net1330),
    .Y(_03034_));
 sky130_fd_sc_hd__o21ai_1 _17892_ (.A1(_03024_),
    .A2(_03033_),
    .B1(net1331),
    .Y(_00231_));
 sky130_fd_sc_hd__a211o_1 _17893_ (.A1(_02938_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03015_),
    .X(_03035_));
 sky130_fd_sc_hd__nand2_1 _17894_ (.A(_03000_),
    .B(net1588),
    .Y(_03036_));
 sky130_fd_sc_hd__o21ai_1 _17895_ (.A1(_03024_),
    .A2(_03035_),
    .B1(net1589),
    .Y(_00232_));
 sky130_fd_sc_hd__a211o_1 _17896_ (.A1(_02943_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03018_),
    .X(_03037_));
 sky130_fd_sc_hd__nand2_1 _17897_ (.A(_03000_),
    .B(net1748),
    .Y(_03038_));
 sky130_fd_sc_hd__o21ai_1 _17898_ (.A1(_03024_),
    .A2(_03037_),
    .B1(net1749),
    .Y(_00233_));
 sky130_fd_sc_hd__a211o_1 _17899_ (.A1(_02948_),
    .A2(_02996_),
    .B1(_03005_),
    .C1(_03021_),
    .X(_03039_));
 sky130_fd_sc_hd__nand2_1 _17900_ (.A(_03000_),
    .B(net1690),
    .Y(_03040_));
 sky130_fd_sc_hd__o21ai_1 _17901_ (.A1(_03024_),
    .A2(_03039_),
    .B1(net1691),
    .Y(_00234_));
 sky130_fd_sc_hd__a211o_1 _17902_ (.A1(_02952_),
    .A2(_02997_),
    .B1(_03005_),
    .C1(_02998_),
    .X(_03041_));
 sky130_fd_sc_hd__nand2_1 _17903_ (.A(_02995_),
    .B(net1850),
    .Y(_03042_));
 sky130_fd_sc_hd__o21ai_1 _17904_ (.A1(_03024_),
    .A2(_03041_),
    .B1(net1851),
    .Y(_00235_));
 sky130_fd_sc_hd__a211o_1 _17905_ (.A1(_02956_),
    .A2(_02997_),
    .B1(_03005_),
    .C1(_03002_),
    .X(_03043_));
 sky130_fd_sc_hd__nand2_1 _17906_ (.A(_02995_),
    .B(net1935),
    .Y(_03044_));
 sky130_fd_sc_hd__o21ai_1 _17907_ (.A1(_03024_),
    .A2(_03043_),
    .B1(net1936),
    .Y(_00236_));
 sky130_fd_sc_hd__buf_4 _17908_ (.A(_09129_),
    .X(_03045_));
 sky130_fd_sc_hd__a211o_1 _17909_ (.A1(_02960_),
    .A2(_02997_),
    .B1(_03045_),
    .C1(_03006_),
    .X(_03046_));
 sky130_fd_sc_hd__nand2_1 _17910_ (.A(_02995_),
    .B(net842),
    .Y(_03047_));
 sky130_fd_sc_hd__o21ai_1 _17911_ (.A1(_03024_),
    .A2(_03046_),
    .B1(net843),
    .Y(_00237_));
 sky130_fd_sc_hd__a211o_1 _17912_ (.A1(_02964_),
    .A2(_02997_),
    .B1(_03045_),
    .C1(_03009_),
    .X(_03048_));
 sky130_fd_sc_hd__nand2_1 _17913_ (.A(_02995_),
    .B(net1852),
    .Y(_03049_));
 sky130_fd_sc_hd__o21ai_1 _17914_ (.A1(_03024_),
    .A2(_03048_),
    .B1(net1853),
    .Y(_00238_));
 sky130_fd_sc_hd__a211o_1 _17915_ (.A1(_02968_),
    .A2(_02997_),
    .B1(_03045_),
    .C1(_03012_),
    .X(_03050_));
 sky130_fd_sc_hd__nand2_1 _17916_ (.A(_02995_),
    .B(net1971),
    .Y(_03051_));
 sky130_fd_sc_hd__o21ai_1 _17917_ (.A1(_03024_),
    .A2(_03050_),
    .B1(_03051_),
    .Y(_00239_));
 sky130_fd_sc_hd__a211o_1 _17918_ (.A1(_02972_),
    .A2(_02997_),
    .B1(_03045_),
    .C1(_03015_),
    .X(_03052_));
 sky130_fd_sc_hd__nand2_1 _17919_ (.A(_02995_),
    .B(net1758),
    .Y(_03053_));
 sky130_fd_sc_hd__o21ai_1 _17920_ (.A1(_03024_),
    .A2(_03052_),
    .B1(net1759),
    .Y(_00240_));
 sky130_fd_sc_hd__a211o_1 _17921_ (.A1(_02976_),
    .A2(_02997_),
    .B1(_03045_),
    .C1(_03018_),
    .X(_03054_));
 sky130_fd_sc_hd__nand2_1 _17922_ (.A(_02995_),
    .B(net1026),
    .Y(_03055_));
 sky130_fd_sc_hd__o21ai_1 _17923_ (.A1(_03024_),
    .A2(_03054_),
    .B1(net1027),
    .Y(_00241_));
 sky130_fd_sc_hd__a211o_1 _17924_ (.A1(_02980_),
    .A2(_02997_),
    .B1(_03045_),
    .C1(_03021_),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _17925_ (.A(_02995_),
    .B(net1040),
    .Y(_03057_));
 sky130_fd_sc_hd__o21ai_1 _17926_ (.A1(_03024_),
    .A2(_03056_),
    .B1(net1041),
    .Y(_00242_));
 sky130_fd_sc_hd__nor2_1 _17927_ (.A(_12292_),
    .B(_02814_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_2 _17928_ (.A(_03058_),
    .B(_09071_),
    .Y(_03059_));
 sky130_fd_sc_hd__inv_2 _17929_ (.A(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__o21ai_4 _17930_ (.A1(_12290_),
    .A2(_03060_),
    .B1(_02818_),
    .Y(_03061_));
 sky130_fd_sc_hd__mux2_1 _17931_ (.A0(_02810_),
    .A1(net2686),
    .S(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _17932_ (.A(_03062_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _17933_ (.A0(_02823_),
    .A1(net2939),
    .S(_03061_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _17934_ (.A(_03063_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _17935_ (.A0(_02827_),
    .A1(net2347),
    .S(_03061_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _17936_ (.A(_03064_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _17937_ (.A0(_02831_),
    .A1(net2676),
    .S(_03061_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _17938_ (.A(_03065_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _17939_ (.A0(_02835_),
    .A1(net2943),
    .S(_03061_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _17940_ (.A(_03066_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _17941_ (.A0(_02839_),
    .A1(net2991),
    .S(_03061_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _17942_ (.A(_03067_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _17943_ (.A0(_02843_),
    .A1(net2374),
    .S(_03061_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _17944_ (.A(_03068_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _17945_ (.A0(_02847_),
    .A1(net2898),
    .S(_03061_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _17946_ (.A(_03069_),
    .X(_00250_));
 sky130_fd_sc_hd__buf_4 _17947_ (.A(_03061_),
    .X(_03070_));
 sky130_fd_sc_hd__buf_4 _17948_ (.A(_03060_),
    .X(_03071_));
 sky130_fd_sc_hd__buf_4 _17949_ (.A(_03060_),
    .X(_03072_));
 sky130_fd_sc_hd__nor2_1 _17950_ (.A(_02854_),
    .B(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__a211o_1 _17951_ (.A1(_02852_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__buf_4 _17952_ (.A(_03061_),
    .X(_03075_));
 sky130_fd_sc_hd__nand2_1 _17953_ (.A(_03075_),
    .B(net1572),
    .Y(_03076_));
 sky130_fd_sc_hd__o21ai_1 _17954_ (.A1(_03070_),
    .A2(_03074_),
    .B1(net1573),
    .Y(_00251_));
 sky130_fd_sc_hd__nor2_1 _17955_ (.A(_02863_),
    .B(_03072_),
    .Y(_03077_));
 sky130_fd_sc_hd__a211o_1 _17956_ (.A1(_02862_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__nand2_1 _17957_ (.A(_03075_),
    .B(net1184),
    .Y(_03079_));
 sky130_fd_sc_hd__o21ai_1 _17958_ (.A1(_03070_),
    .A2(_03078_),
    .B1(net1185),
    .Y(_00252_));
 sky130_fd_sc_hd__nor2_1 _17959_ (.A(_02870_),
    .B(_03072_),
    .Y(_03080_));
 sky130_fd_sc_hd__a211o_1 _17960_ (.A1(_02869_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__nand2_1 _17961_ (.A(_03075_),
    .B(net1530),
    .Y(_03082_));
 sky130_fd_sc_hd__o21ai_1 _17962_ (.A1(_03070_),
    .A2(_03081_),
    .B1(net1531),
    .Y(_00253_));
 sky130_fd_sc_hd__nor2_1 _17963_ (.A(_02877_),
    .B(_03072_),
    .Y(_03083_));
 sky130_fd_sc_hd__a211o_1 _17964_ (.A1(_02876_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__nand2_1 _17965_ (.A(_03075_),
    .B(net830),
    .Y(_03085_));
 sky130_fd_sc_hd__o21ai_1 _17966_ (.A1(_03070_),
    .A2(_03084_),
    .B1(net831),
    .Y(_00254_));
 sky130_fd_sc_hd__nor2_1 _17967_ (.A(_02884_),
    .B(_03072_),
    .Y(_03086_));
 sky130_fd_sc_hd__a211o_1 _17968_ (.A1(_02883_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__nand2_1 _17969_ (.A(_03075_),
    .B(net1264),
    .Y(_03088_));
 sky130_fd_sc_hd__o21ai_1 _17970_ (.A1(_03070_),
    .A2(_03087_),
    .B1(net1265),
    .Y(_00255_));
 sky130_fd_sc_hd__nor2_1 _17971_ (.A(_02891_),
    .B(_03072_),
    .Y(_03089_));
 sky130_fd_sc_hd__a211o_1 _17972_ (.A1(_02890_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__nand2_1 _17973_ (.A(_03075_),
    .B(net1018),
    .Y(_03091_));
 sky130_fd_sc_hd__o21ai_1 _17974_ (.A1(_03070_),
    .A2(_03090_),
    .B1(net1019),
    .Y(_00256_));
 sky130_fd_sc_hd__nor2_1 _17975_ (.A(_02898_),
    .B(_03072_),
    .Y(_03092_));
 sky130_fd_sc_hd__a211o_1 _17976_ (.A1(_02897_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__nand2_1 _17977_ (.A(_03075_),
    .B(net1512),
    .Y(_03094_));
 sky130_fd_sc_hd__o21ai_1 _17978_ (.A1(_03070_),
    .A2(_03093_),
    .B1(net1513),
    .Y(_00257_));
 sky130_fd_sc_hd__nor2_1 _17979_ (.A(_02905_),
    .B(_03072_),
    .Y(_03095_));
 sky130_fd_sc_hd__a211o_1 _17980_ (.A1(_02904_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__nand2_1 _17981_ (.A(_03075_),
    .B(net1682),
    .Y(_03097_));
 sky130_fd_sc_hd__o21ai_1 _17982_ (.A1(_03070_),
    .A2(_03096_),
    .B1(net1683),
    .Y(_00258_));
 sky130_fd_sc_hd__buf_4 _17983_ (.A(_03061_),
    .X(_03098_));
 sky130_fd_sc_hd__a211o_1 _17984_ (.A1(_02912_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03073_),
    .X(_03099_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(_03075_),
    .B(net780),
    .Y(_03100_));
 sky130_fd_sc_hd__o21ai_1 _17986_ (.A1(_03098_),
    .A2(_03099_),
    .B1(net781),
    .Y(_00259_));
 sky130_fd_sc_hd__a211o_1 _17987_ (.A1(_02917_),
    .A2(_03071_),
    .B1(_03045_),
    .C1(_03077_),
    .X(_03101_));
 sky130_fd_sc_hd__nand2_1 _17988_ (.A(_03075_),
    .B(net596),
    .Y(_03102_));
 sky130_fd_sc_hd__o21ai_1 _17989_ (.A1(_03098_),
    .A2(_03101_),
    .B1(net597),
    .Y(_00260_));
 sky130_fd_sc_hd__buf_4 _17990_ (.A(_09129_),
    .X(_03103_));
 sky130_fd_sc_hd__a211o_1 _17991_ (.A1(_02922_),
    .A2(_03071_),
    .B1(_03103_),
    .C1(_03080_),
    .X(_03104_));
 sky130_fd_sc_hd__nand2_1 _17992_ (.A(_03075_),
    .B(net646),
    .Y(_03105_));
 sky130_fd_sc_hd__o21ai_1 _17993_ (.A1(_03098_),
    .A2(_03104_),
    .B1(net647),
    .Y(_00261_));
 sky130_fd_sc_hd__a211o_1 _17994_ (.A1(_02928_),
    .A2(_03071_),
    .B1(_03103_),
    .C1(_03083_),
    .X(_03106_));
 sky130_fd_sc_hd__nand2_1 _17995_ (.A(_03075_),
    .B(net810),
    .Y(_03107_));
 sky130_fd_sc_hd__o21ai_1 _17996_ (.A1(_03098_),
    .A2(_03106_),
    .B1(net811),
    .Y(_00262_));
 sky130_fd_sc_hd__a211o_1 _17997_ (.A1(_02933_),
    .A2(_03071_),
    .B1(_03103_),
    .C1(_03086_),
    .X(_03108_));
 sky130_fd_sc_hd__nand2_1 _17998_ (.A(_03075_),
    .B(net1170),
    .Y(_03109_));
 sky130_fd_sc_hd__o21ai_1 _17999_ (.A1(_03098_),
    .A2(_03108_),
    .B1(net1171),
    .Y(_00263_));
 sky130_fd_sc_hd__a211o_1 _18000_ (.A1(_02938_),
    .A2(_03071_),
    .B1(_03103_),
    .C1(_03089_),
    .X(_03110_));
 sky130_fd_sc_hd__nand2_1 _18001_ (.A(_03075_),
    .B(net818),
    .Y(_03111_));
 sky130_fd_sc_hd__o21ai_1 _18002_ (.A1(_03098_),
    .A2(_03110_),
    .B1(net819),
    .Y(_00264_));
 sky130_fd_sc_hd__a211o_1 _18003_ (.A1(_02943_),
    .A2(_03071_),
    .B1(_03103_),
    .C1(_03092_),
    .X(_03112_));
 sky130_fd_sc_hd__nand2_1 _18004_ (.A(_03075_),
    .B(net1883),
    .Y(_03113_));
 sky130_fd_sc_hd__o21ai_1 _18005_ (.A1(_03098_),
    .A2(_03112_),
    .B1(net1884),
    .Y(_00265_));
 sky130_fd_sc_hd__a211o_1 _18006_ (.A1(_02948_),
    .A2(_03071_),
    .B1(_03103_),
    .C1(_03095_),
    .X(_03114_));
 sky130_fd_sc_hd__nand2_1 _18007_ (.A(_03075_),
    .B(net840),
    .Y(_03115_));
 sky130_fd_sc_hd__o21ai_1 _18008_ (.A1(_03098_),
    .A2(_03114_),
    .B1(net841),
    .Y(_00266_));
 sky130_fd_sc_hd__a211o_1 _18009_ (.A1(_02952_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03073_),
    .X(_03116_));
 sky130_fd_sc_hd__nand2_1 _18010_ (.A(_03070_),
    .B(net640),
    .Y(_03117_));
 sky130_fd_sc_hd__o21ai_1 _18011_ (.A1(_03098_),
    .A2(_03116_),
    .B1(net641),
    .Y(_00267_));
 sky130_fd_sc_hd__a211o_1 _18012_ (.A1(_02956_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03077_),
    .X(_03118_));
 sky130_fd_sc_hd__nand2_1 _18013_ (.A(_03070_),
    .B(net584),
    .Y(_03119_));
 sky130_fd_sc_hd__o21ai_1 _18014_ (.A1(_03098_),
    .A2(_03118_),
    .B1(net585),
    .Y(_00268_));
 sky130_fd_sc_hd__a211o_1 _18015_ (.A1(_02960_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03080_),
    .X(_03120_));
 sky130_fd_sc_hd__nand2_1 _18016_ (.A(_03070_),
    .B(net624),
    .Y(_03121_));
 sky130_fd_sc_hd__o21ai_1 _18017_ (.A1(_03098_),
    .A2(_03120_),
    .B1(net625),
    .Y(_00269_));
 sky130_fd_sc_hd__a211o_1 _18018_ (.A1(_02964_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03083_),
    .X(_03122_));
 sky130_fd_sc_hd__nand2_1 _18019_ (.A(_03070_),
    .B(net1937),
    .Y(_03123_));
 sky130_fd_sc_hd__o21ai_1 _18020_ (.A1(_03098_),
    .A2(_03122_),
    .B1(net1938),
    .Y(_00270_));
 sky130_fd_sc_hd__a211o_1 _18021_ (.A1(_02968_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03086_),
    .X(_03124_));
 sky130_fd_sc_hd__nand2_1 _18022_ (.A(_03070_),
    .B(net1895),
    .Y(_03125_));
 sky130_fd_sc_hd__o21ai_1 _18023_ (.A1(_03098_),
    .A2(_03124_),
    .B1(net1896),
    .Y(_00271_));
 sky130_fd_sc_hd__a211o_1 _18024_ (.A1(_02972_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03089_),
    .X(_03126_));
 sky130_fd_sc_hd__nand2_1 _18025_ (.A(_03070_),
    .B(net550),
    .Y(_03127_));
 sky130_fd_sc_hd__o21ai_1 _18026_ (.A1(_03098_),
    .A2(_03126_),
    .B1(net551),
    .Y(_00272_));
 sky130_fd_sc_hd__a211o_1 _18027_ (.A1(_02976_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03092_),
    .X(_03128_));
 sky130_fd_sc_hd__nand2_1 _18028_ (.A(_03070_),
    .B(net1502),
    .Y(_03129_));
 sky130_fd_sc_hd__o21ai_1 _18029_ (.A1(_03098_),
    .A2(_03128_),
    .B1(net1503),
    .Y(_00273_));
 sky130_fd_sc_hd__a211o_1 _18030_ (.A1(_02980_),
    .A2(_03072_),
    .B1(_03103_),
    .C1(_03095_),
    .X(_03130_));
 sky130_fd_sc_hd__nand2_1 _18031_ (.A(_03070_),
    .B(net730),
    .Y(_03131_));
 sky130_fd_sc_hd__o21ai_1 _18032_ (.A1(_03098_),
    .A2(_03130_),
    .B1(net731),
    .Y(_00274_));
 sky130_fd_sc_hd__nor2_1 _18033_ (.A(_12171_),
    .B(_02814_),
    .Y(_03132_));
 sky130_fd_sc_hd__inv_2 _18034_ (.A(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__nor2_4 _18035_ (.A(_12177_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__o21ai_4 _18036_ (.A1(_12290_),
    .A2(_03134_),
    .B1(_02818_),
    .Y(_03135_));
 sky130_fd_sc_hd__mux2_1 _18037_ (.A0(_02810_),
    .A1(net2713),
    .S(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_1 _18038_ (.A(_03136_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _18039_ (.A0(_02823_),
    .A1(net2190),
    .S(_03135_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_1 _18040_ (.A(_03137_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _18041_ (.A0(_02827_),
    .A1(net2317),
    .S(_03135_),
    .X(_03138_));
 sky130_fd_sc_hd__clkbuf_1 _18042_ (.A(_03138_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _18043_ (.A0(_02831_),
    .A1(net2322),
    .S(_03135_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_1 _18044_ (.A(_03139_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _18045_ (.A0(_02835_),
    .A1(net2222),
    .S(_03135_),
    .X(_03140_));
 sky130_fd_sc_hd__clkbuf_1 _18046_ (.A(_03140_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _18047_ (.A0(_02839_),
    .A1(net2157),
    .S(_03135_),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_1 _18048_ (.A(_03141_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _18049_ (.A0(_02843_),
    .A1(net3198),
    .S(_03135_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_1 _18050_ (.A(_03142_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _18051_ (.A0(_02847_),
    .A1(net2105),
    .S(_03135_),
    .X(_03143_));
 sky130_fd_sc_hd__clkbuf_1 _18052_ (.A(_03143_),
    .X(_00282_));
 sky130_fd_sc_hd__buf_4 _18053_ (.A(_03135_),
    .X(_03144_));
 sky130_fd_sc_hd__buf_4 _18054_ (.A(_03134_),
    .X(_03145_));
 sky130_fd_sc_hd__buf_4 _18055_ (.A(_03134_),
    .X(_03146_));
 sky130_fd_sc_hd__nor2_1 _18056_ (.A(_02854_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__a211o_1 _18057_ (.A1(_02852_),
    .A2(_03145_),
    .B1(_03103_),
    .C1(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__buf_4 _18058_ (.A(_03135_),
    .X(_03149_));
 sky130_fd_sc_hd__nand2_1 _18059_ (.A(_03149_),
    .B(net1897),
    .Y(_03150_));
 sky130_fd_sc_hd__o21ai_1 _18060_ (.A1(_03144_),
    .A2(_03148_),
    .B1(net1898),
    .Y(_00283_));
 sky130_fd_sc_hd__nor2_1 _18061_ (.A(_02863_),
    .B(_03146_),
    .Y(_03151_));
 sky130_fd_sc_hd__a211o_1 _18062_ (.A1(_02862_),
    .A2(_03145_),
    .B1(_03103_),
    .C1(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__nand2_1 _18063_ (.A(_03149_),
    .B(net1911),
    .Y(_03153_));
 sky130_fd_sc_hd__o21ai_1 _18064_ (.A1(_03144_),
    .A2(_03152_),
    .B1(net1912),
    .Y(_00284_));
 sky130_fd_sc_hd__buf_4 _18065_ (.A(_09129_),
    .X(_03154_));
 sky130_fd_sc_hd__nor2_1 _18066_ (.A(_02870_),
    .B(_03146_),
    .Y(_03155_));
 sky130_fd_sc_hd__a211o_1 _18067_ (.A1(_02869_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__nand2_1 _18068_ (.A(_03149_),
    .B(net1955),
    .Y(_03157_));
 sky130_fd_sc_hd__o21ai_1 _18069_ (.A1(_03144_),
    .A2(_03156_),
    .B1(_03157_),
    .Y(_00285_));
 sky130_fd_sc_hd__nor2_1 _18070_ (.A(_02877_),
    .B(_03146_),
    .Y(_03158_));
 sky130_fd_sc_hd__a211o_1 _18071_ (.A1(_02876_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__nand2_1 _18072_ (.A(_03149_),
    .B(net1550),
    .Y(_03160_));
 sky130_fd_sc_hd__o21ai_1 _18073_ (.A1(_03144_),
    .A2(_03159_),
    .B1(net1551),
    .Y(_00286_));
 sky130_fd_sc_hd__nor2_1 _18074_ (.A(_02884_),
    .B(_03146_),
    .Y(_03161_));
 sky130_fd_sc_hd__a211o_1 _18075_ (.A1(_02883_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__nand2_1 _18076_ (.A(_03149_),
    .B(net1292),
    .Y(_03163_));
 sky130_fd_sc_hd__o21ai_1 _18077_ (.A1(_03144_),
    .A2(_03162_),
    .B1(net1293),
    .Y(_00287_));
 sky130_fd_sc_hd__nor2_1 _18078_ (.A(_02891_),
    .B(_03146_),
    .Y(_03164_));
 sky130_fd_sc_hd__a211o_1 _18079_ (.A1(_02890_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__nand2_1 _18080_ (.A(_03149_),
    .B(net1983),
    .Y(_03166_));
 sky130_fd_sc_hd__o21ai_1 _18081_ (.A1(_03144_),
    .A2(_03165_),
    .B1(_03166_),
    .Y(_00288_));
 sky130_fd_sc_hd__nor2_1 _18082_ (.A(_02898_),
    .B(_03146_),
    .Y(_03167_));
 sky130_fd_sc_hd__a211o_1 _18083_ (.A1(_02897_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__nand2_1 _18084_ (.A(_03149_),
    .B(net1158),
    .Y(_03169_));
 sky130_fd_sc_hd__o21ai_1 _18085_ (.A1(_03144_),
    .A2(_03168_),
    .B1(net1159),
    .Y(_00289_));
 sky130_fd_sc_hd__nor2_1 _18086_ (.A(_02905_),
    .B(_03146_),
    .Y(_03170_));
 sky130_fd_sc_hd__a211o_1 _18087_ (.A1(_02904_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__nand2_1 _18088_ (.A(_03149_),
    .B(net1974),
    .Y(_03172_));
 sky130_fd_sc_hd__o21ai_1 _18089_ (.A1(_03144_),
    .A2(_03171_),
    .B1(_03172_),
    .Y(_00290_));
 sky130_fd_sc_hd__buf_4 _18090_ (.A(_03135_),
    .X(_03173_));
 sky130_fd_sc_hd__a211o_1 _18091_ (.A1(_02912_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03147_),
    .X(_03174_));
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(_03149_),
    .B(net1968),
    .Y(_03175_));
 sky130_fd_sc_hd__o21ai_1 _18093_ (.A1(_03173_),
    .A2(_03174_),
    .B1(_03175_),
    .Y(_00291_));
 sky130_fd_sc_hd__a211o_1 _18094_ (.A1(_02917_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03151_),
    .X(_03176_));
 sky130_fd_sc_hd__nand2_1 _18095_ (.A(_03149_),
    .B(net1970),
    .Y(_03177_));
 sky130_fd_sc_hd__o21ai_1 _18096_ (.A1(_03173_),
    .A2(_03176_),
    .B1(_03177_),
    .Y(_00292_));
 sky130_fd_sc_hd__a211o_1 _18097_ (.A1(_02922_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03155_),
    .X(_03178_));
 sky130_fd_sc_hd__nand2_1 _18098_ (.A(_03149_),
    .B(net1976),
    .Y(_03179_));
 sky130_fd_sc_hd__o21ai_1 _18099_ (.A1(_03173_),
    .A2(_03178_),
    .B1(_03179_),
    .Y(_00293_));
 sky130_fd_sc_hd__a211o_1 _18100_ (.A1(_02928_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03158_),
    .X(_03180_));
 sky130_fd_sc_hd__nand2_1 _18101_ (.A(_03149_),
    .B(net1742),
    .Y(_03181_));
 sky130_fd_sc_hd__o21ai_1 _18102_ (.A1(_03173_),
    .A2(_03180_),
    .B1(net1743),
    .Y(_00294_));
 sky130_fd_sc_hd__a211o_1 _18103_ (.A1(_02933_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03161_),
    .X(_03182_));
 sky130_fd_sc_hd__nand2_1 _18104_ (.A(_03149_),
    .B(net912),
    .Y(_03183_));
 sky130_fd_sc_hd__o21ai_1 _18105_ (.A1(_03173_),
    .A2(_03182_),
    .B1(net913),
    .Y(_00295_));
 sky130_fd_sc_hd__a211o_1 _18106_ (.A1(_02938_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03164_),
    .X(_03184_));
 sky130_fd_sc_hd__nand2_1 _18107_ (.A(_03149_),
    .B(net1982),
    .Y(_03185_));
 sky130_fd_sc_hd__o21ai_1 _18108_ (.A1(_03173_),
    .A2(_03184_),
    .B1(_03185_),
    .Y(_00296_));
 sky130_fd_sc_hd__a211o_1 _18109_ (.A1(_02943_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03167_),
    .X(_03186_));
 sky130_fd_sc_hd__nand2_1 _18110_ (.A(_03149_),
    .B(net1542),
    .Y(_03187_));
 sky130_fd_sc_hd__o21ai_1 _18111_ (.A1(_03173_),
    .A2(_03186_),
    .B1(net1543),
    .Y(_00297_));
 sky130_fd_sc_hd__a211o_1 _18112_ (.A1(_02948_),
    .A2(_03145_),
    .B1(_03154_),
    .C1(_03170_),
    .X(_03188_));
 sky130_fd_sc_hd__nand2_1 _18113_ (.A(_03149_),
    .B(net1990),
    .Y(_03189_));
 sky130_fd_sc_hd__o21ai_1 _18114_ (.A1(_03173_),
    .A2(_03188_),
    .B1(_03189_),
    .Y(_00298_));
 sky130_fd_sc_hd__a211o_1 _18115_ (.A1(_02952_),
    .A2(_03146_),
    .B1(_03154_),
    .C1(_03147_),
    .X(_03190_));
 sky130_fd_sc_hd__nand2_1 _18116_ (.A(_03144_),
    .B(net1975),
    .Y(_03191_));
 sky130_fd_sc_hd__o21ai_1 _18117_ (.A1(_03173_),
    .A2(_03190_),
    .B1(_03191_),
    .Y(_00299_));
 sky130_fd_sc_hd__a211o_1 _18118_ (.A1(_02956_),
    .A2(_03146_),
    .B1(_03154_),
    .C1(_03151_),
    .X(_03192_));
 sky130_fd_sc_hd__nand2_1 _18119_ (.A(_03144_),
    .B(net1981),
    .Y(_03193_));
 sky130_fd_sc_hd__o21ai_1 _18120_ (.A1(_03173_),
    .A2(_03192_),
    .B1(_03193_),
    .Y(_00300_));
 sky130_fd_sc_hd__clkbuf_8 _18121_ (.A(_09129_),
    .X(_03194_));
 sky130_fd_sc_hd__a211o_1 _18122_ (.A1(_02960_),
    .A2(_03146_),
    .B1(_03194_),
    .C1(_03155_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2_1 _18123_ (.A(_03144_),
    .B(net1984),
    .Y(_03196_));
 sky130_fd_sc_hd__o21ai_1 _18124_ (.A1(_03173_),
    .A2(_03195_),
    .B1(_03196_),
    .Y(_00301_));
 sky130_fd_sc_hd__a211o_1 _18125_ (.A1(_02964_),
    .A2(_03146_),
    .B1(_03194_),
    .C1(_03158_),
    .X(_03197_));
 sky130_fd_sc_hd__nand2_1 _18126_ (.A(_03144_),
    .B(net1944),
    .Y(_03198_));
 sky130_fd_sc_hd__o21ai_1 _18127_ (.A1(_03173_),
    .A2(_03197_),
    .B1(net1945),
    .Y(_00302_));
 sky130_fd_sc_hd__a211o_1 _18128_ (.A1(_02968_),
    .A2(_03146_),
    .B1(_03194_),
    .C1(_03161_),
    .X(_03199_));
 sky130_fd_sc_hd__nand2_1 _18129_ (.A(_03144_),
    .B(net1887),
    .Y(_03200_));
 sky130_fd_sc_hd__o21ai_1 _18130_ (.A1(_03173_),
    .A2(_03199_),
    .B1(net1888),
    .Y(_00303_));
 sky130_fd_sc_hd__a211o_1 _18131_ (.A1(_02972_),
    .A2(_03146_),
    .B1(_03194_),
    .C1(_03164_),
    .X(_03201_));
 sky130_fd_sc_hd__nand2_1 _18132_ (.A(_03144_),
    .B(net1582),
    .Y(_03202_));
 sky130_fd_sc_hd__o21ai_1 _18133_ (.A1(_03173_),
    .A2(_03201_),
    .B1(net1583),
    .Y(_00304_));
 sky130_fd_sc_hd__a211o_1 _18134_ (.A1(_02976_),
    .A2(_03146_),
    .B1(_03194_),
    .C1(_03167_),
    .X(_03203_));
 sky130_fd_sc_hd__nand2_1 _18135_ (.A(_03144_),
    .B(net1304),
    .Y(_03204_));
 sky130_fd_sc_hd__o21ai_1 _18136_ (.A1(_03173_),
    .A2(_03203_),
    .B1(net1305),
    .Y(_00305_));
 sky130_fd_sc_hd__a211o_1 _18137_ (.A1(_02980_),
    .A2(_03146_),
    .B1(_03194_),
    .C1(_03170_),
    .X(_03205_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(_03144_),
    .B(net1907),
    .Y(_03206_));
 sky130_fd_sc_hd__o21ai_1 _18139_ (.A1(_03173_),
    .A2(_03205_),
    .B1(net1908),
    .Y(_00306_));
 sky130_fd_sc_hd__nor2_2 _18140_ (.A(\line_cache_idx[5] ),
    .B(_09090_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_1 _18141_ (.A(_03207_),
    .B(_12174_),
    .Y(_03208_));
 sky130_fd_sc_hd__or2_1 _18142_ (.A(_02812_),
    .B(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__inv_2 _18143_ (.A(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_2 _18144_ (.A(_03210_),
    .B(_12313_),
    .Y(_03211_));
 sky130_fd_sc_hd__a21bo_1 _18145_ (.A1(_03211_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_8 _18146_ (.A(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_1 _18147_ (.A0(_02810_),
    .A1(net3580),
    .S(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_1 _18148_ (.A(_03214_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _18149_ (.A0(_02823_),
    .A1(net2241),
    .S(_03213_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _18150_ (.A(_03215_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _18151_ (.A0(_02827_),
    .A1(net2417),
    .S(_03213_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_1 _18152_ (.A(_03216_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _18153_ (.A0(_02831_),
    .A1(net2763),
    .S(_03213_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_1 _18154_ (.A(_03217_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _18155_ (.A0(_02835_),
    .A1(net3373),
    .S(_03213_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_1 _18156_ (.A(_03218_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _18157_ (.A0(_02839_),
    .A1(net3697),
    .S(_03213_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_1 _18158_ (.A(_03219_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _18159_ (.A0(_02843_),
    .A1(net2733),
    .S(_03213_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_1 _18160_ (.A(_03220_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _18161_ (.A0(_02847_),
    .A1(net2677),
    .S(_03213_),
    .X(_03221_));
 sky130_fd_sc_hd__clkbuf_1 _18162_ (.A(_03221_),
    .X(_00314_));
 sky130_fd_sc_hd__clkbuf_16 _18163_ (.A(_02850_),
    .X(_03222_));
 sky130_fd_sc_hd__buf_4 _18164_ (.A(_03211_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_4 _18165_ (.A(_03211_),
    .X(_03224_));
 sky130_fd_sc_hd__nand2_1 _18166_ (.A(_03224_),
    .B(_12185_),
    .Y(_03225_));
 sky130_fd_sc_hd__o211a_1 _18167_ (.A1(_03222_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _18168_ (.A0(_03226_),
    .A1(net3469),
    .S(_03213_),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_1 _18169_ (.A(_03227_),
    .X(_00315_));
 sky130_fd_sc_hd__clkbuf_16 _18170_ (.A(_02860_),
    .X(_03228_));
 sky130_fd_sc_hd__nand2_1 _18171_ (.A(_03224_),
    .B(_12198_),
    .Y(_03229_));
 sky130_fd_sc_hd__o211a_1 _18172_ (.A1(_03228_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _18173_ (.A0(_03230_),
    .A1(net3572),
    .S(_03213_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_1 _18174_ (.A(_03231_),
    .X(_00316_));
 sky130_fd_sc_hd__buf_12 _18175_ (.A(_02867_),
    .X(_03232_));
 sky130_fd_sc_hd__nand2_1 _18176_ (.A(_03224_),
    .B(_12206_),
    .Y(_03233_));
 sky130_fd_sc_hd__o211a_1 _18177_ (.A1(_03232_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _18178_ (.A0(_03234_),
    .A1(net3273),
    .S(_03213_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_1 _18179_ (.A(_03235_),
    .X(_00317_));
 sky130_fd_sc_hd__buf_12 _18180_ (.A(_02874_),
    .X(_03236_));
 sky130_fd_sc_hd__nand2_1 _18181_ (.A(_03224_),
    .B(_12214_),
    .Y(_03237_));
 sky130_fd_sc_hd__o211a_1 _18182_ (.A1(_03236_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _18183_ (.A0(_03238_),
    .A1(net3501),
    .S(_03213_),
    .X(_03239_));
 sky130_fd_sc_hd__clkbuf_1 _18184_ (.A(_03239_),
    .X(_00318_));
 sky130_fd_sc_hd__clkbuf_16 _18185_ (.A(_02881_),
    .X(_03240_));
 sky130_fd_sc_hd__nand2_1 _18186_ (.A(_03224_),
    .B(_12222_),
    .Y(_03241_));
 sky130_fd_sc_hd__o211a_1 _18187_ (.A1(_03240_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__mux2_1 _18188_ (.A0(_03242_),
    .A1(net3512),
    .S(_03213_),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_1 _18189_ (.A(_03243_),
    .X(_00319_));
 sky130_fd_sc_hd__buf_12 _18190_ (.A(_02888_),
    .X(_03244_));
 sky130_fd_sc_hd__nand2_1 _18191_ (.A(_03224_),
    .B(_12230_),
    .Y(_03245_));
 sky130_fd_sc_hd__o211a_1 _18192_ (.A1(_03244_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _18193_ (.A0(_03246_),
    .A1(net2474),
    .S(_03213_),
    .X(_03247_));
 sky130_fd_sc_hd__clkbuf_1 _18194_ (.A(_03247_),
    .X(_00320_));
 sky130_fd_sc_hd__buf_12 _18195_ (.A(_02895_),
    .X(_03248_));
 sky130_fd_sc_hd__nand2_1 _18196_ (.A(_03224_),
    .B(_12238_),
    .Y(_03249_));
 sky130_fd_sc_hd__o211a_1 _18197_ (.A1(_03248_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_1 _18198_ (.A0(_03250_),
    .A1(net2693),
    .S(_03213_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_1 _18199_ (.A(_03251_),
    .X(_00321_));
 sky130_fd_sc_hd__clkbuf_16 _18200_ (.A(_02902_),
    .X(_03252_));
 sky130_fd_sc_hd__nand2_1 _18201_ (.A(_03224_),
    .B(_12246_),
    .Y(_03253_));
 sky130_fd_sc_hd__o211a_1 _18202_ (.A1(_03252_),
    .A2(_03223_),
    .B1(_12181_),
    .C1(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _18203_ (.A0(_03254_),
    .A1(net3027),
    .S(_03213_),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_1 _18204_ (.A(_03255_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_12 _18205_ (.A(_02910_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_4 _18206_ (.A(_12180_),
    .X(_03257_));
 sky130_fd_sc_hd__o211a_1 _18207_ (.A1(_03256_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03225_),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_8 _18208_ (.A(_03212_),
    .X(_03259_));
 sky130_fd_sc_hd__mux2_1 _18209_ (.A0(_03258_),
    .A1(net2754),
    .S(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__clkbuf_1 _18210_ (.A(_03260_),
    .X(_00323_));
 sky130_fd_sc_hd__clkbuf_16 _18211_ (.A(_02915_),
    .X(_03261_));
 sky130_fd_sc_hd__o211a_1 _18212_ (.A1(_03261_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03229_),
    .X(_03262_));
 sky130_fd_sc_hd__mux2_1 _18213_ (.A0(_03262_),
    .A1(net3212),
    .S(_03259_),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_1 _18214_ (.A(_03263_),
    .X(_00324_));
 sky130_fd_sc_hd__buf_12 _18215_ (.A(_02920_),
    .X(_03264_));
 sky130_fd_sc_hd__o211a_1 _18216_ (.A1(_03264_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03233_),
    .X(_03265_));
 sky130_fd_sc_hd__mux2_1 _18217_ (.A0(_03265_),
    .A1(net3331),
    .S(_03259_),
    .X(_03266_));
 sky130_fd_sc_hd__clkbuf_1 _18218_ (.A(_03266_),
    .X(_00325_));
 sky130_fd_sc_hd__clkbuf_16 _18219_ (.A(_02926_),
    .X(_03267_));
 sky130_fd_sc_hd__o211a_1 _18220_ (.A1(_03267_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03237_),
    .X(_03268_));
 sky130_fd_sc_hd__mux2_1 _18221_ (.A0(_03268_),
    .A1(net2351),
    .S(_03259_),
    .X(_03269_));
 sky130_fd_sc_hd__clkbuf_1 _18222_ (.A(_03269_),
    .X(_00326_));
 sky130_fd_sc_hd__clkbuf_16 _18223_ (.A(_02931_),
    .X(_03270_));
 sky130_fd_sc_hd__o211a_1 _18224_ (.A1(_03270_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03241_),
    .X(_03271_));
 sky130_fd_sc_hd__mux2_1 _18225_ (.A0(_03271_),
    .A1(net2649),
    .S(_03259_),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_1 _18226_ (.A(_03272_),
    .X(_00327_));
 sky130_fd_sc_hd__clkbuf_16 _18227_ (.A(_02936_),
    .X(_03273_));
 sky130_fd_sc_hd__o211a_1 _18228_ (.A1(_03273_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03245_),
    .X(_03274_));
 sky130_fd_sc_hd__mux2_1 _18229_ (.A0(_03274_),
    .A1(net2776),
    .S(_03259_),
    .X(_03275_));
 sky130_fd_sc_hd__clkbuf_1 _18230_ (.A(_03275_),
    .X(_00328_));
 sky130_fd_sc_hd__buf_12 _18231_ (.A(_02941_),
    .X(_03276_));
 sky130_fd_sc_hd__o211a_1 _18232_ (.A1(_03276_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03249_),
    .X(_03277_));
 sky130_fd_sc_hd__mux2_1 _18233_ (.A0(_03277_),
    .A1(net3089),
    .S(_03259_),
    .X(_03278_));
 sky130_fd_sc_hd__clkbuf_1 _18234_ (.A(_03278_),
    .X(_00329_));
 sky130_fd_sc_hd__clkbuf_16 _18235_ (.A(_02946_),
    .X(_03279_));
 sky130_fd_sc_hd__o211a_1 _18236_ (.A1(_03279_),
    .A2(_03223_),
    .B1(_03257_),
    .C1(_03253_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _18237_ (.A0(_03280_),
    .A1(net2501),
    .S(_03259_),
    .X(_03281_));
 sky130_fd_sc_hd__clkbuf_1 _18238_ (.A(_03281_),
    .X(_00330_));
 sky130_fd_sc_hd__o211a_1 _18239_ (.A1(_12170_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03225_),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_1 _18240_ (.A0(_03282_),
    .A1(net2921),
    .S(_03259_),
    .X(_03283_));
 sky130_fd_sc_hd__clkbuf_1 _18241_ (.A(_03283_),
    .X(_00331_));
 sky130_fd_sc_hd__o211a_1 _18242_ (.A1(_12195_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03229_),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _18243_ (.A0(_03284_),
    .A1(net2606),
    .S(_03259_),
    .X(_03285_));
 sky130_fd_sc_hd__clkbuf_1 _18244_ (.A(_03285_),
    .X(_00332_));
 sky130_fd_sc_hd__o211a_1 _18245_ (.A1(_12203_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03233_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _18246_ (.A0(_03286_),
    .A1(net2209),
    .S(_03259_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_1 _18247_ (.A(_03287_),
    .X(_00333_));
 sky130_fd_sc_hd__o211a_1 _18248_ (.A1(_12211_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03237_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _18249_ (.A0(_03288_),
    .A1(net2611),
    .S(_03259_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_1 _18250_ (.A(_03289_),
    .X(_00334_));
 sky130_fd_sc_hd__o211a_1 _18251_ (.A1(_12219_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03241_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _18252_ (.A0(_03290_),
    .A1(net2775),
    .S(_03259_),
    .X(_03291_));
 sky130_fd_sc_hd__clkbuf_1 _18253_ (.A(_03291_),
    .X(_00335_));
 sky130_fd_sc_hd__o211a_1 _18254_ (.A1(_12227_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03245_),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _18255_ (.A0(_03292_),
    .A1(net3317),
    .S(_03259_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_1 _18256_ (.A(_03293_),
    .X(_00336_));
 sky130_fd_sc_hd__o211a_1 _18257_ (.A1(_12235_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03249_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _18258_ (.A0(_03294_),
    .A1(net3183),
    .S(_03259_),
    .X(_03295_));
 sky130_fd_sc_hd__clkbuf_1 _18259_ (.A(_03295_),
    .X(_00337_));
 sky130_fd_sc_hd__o211a_1 _18260_ (.A1(_12243_),
    .A2(_03224_),
    .B1(_03257_),
    .C1(_03253_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _18261_ (.A0(_03296_),
    .A1(net2842),
    .S(_03259_),
    .X(_03297_));
 sky130_fd_sc_hd__clkbuf_1 _18262_ (.A(_03297_),
    .X(_00338_));
 sky130_fd_sc_hd__nor2_1 _18263_ (.A(_12293_),
    .B(_03208_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_2 _18264_ (.A(_03298_),
    .B(_12313_),
    .Y(_03299_));
 sky130_fd_sc_hd__a21bo_1 _18265_ (.A1(_03299_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03300_));
 sky130_fd_sc_hd__clkbuf_8 _18266_ (.A(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _18267_ (.A0(_02810_),
    .A1(net3444),
    .S(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_1 _18268_ (.A(_03302_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _18269_ (.A0(_02823_),
    .A1(net3389),
    .S(_03301_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _18270_ (.A(_03303_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _18271_ (.A0(_02827_),
    .A1(net2433),
    .S(_03301_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _18272_ (.A(_03304_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _18273_ (.A0(_02831_),
    .A1(net3268),
    .S(_03301_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_1 _18274_ (.A(_03305_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _18275_ (.A0(_02835_),
    .A1(net3004),
    .S(_03301_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _18276_ (.A(_03306_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _18277_ (.A0(_02839_),
    .A1(net3400),
    .S(_03301_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _18278_ (.A(_03307_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _18279_ (.A0(_02843_),
    .A1(net3049),
    .S(_03301_),
    .X(_03308_));
 sky130_fd_sc_hd__clkbuf_1 _18280_ (.A(_03308_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(_02847_),
    .A1(net3271),
    .S(_03301_),
    .X(_03309_));
 sky130_fd_sc_hd__clkbuf_1 _18282_ (.A(_03309_),
    .X(_00346_));
 sky130_fd_sc_hd__buf_4 _18283_ (.A(_03299_),
    .X(_03310_));
 sky130_fd_sc_hd__buf_4 _18284_ (.A(_12180_),
    .X(_03311_));
 sky130_fd_sc_hd__buf_4 _18285_ (.A(_03299_),
    .X(_03312_));
 sky130_fd_sc_hd__nand2_1 _18286_ (.A(_03312_),
    .B(_12185_),
    .Y(_03313_));
 sky130_fd_sc_hd__o211a_1 _18287_ (.A1(_03222_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _18288_ (.A0(_03314_),
    .A1(net2361),
    .S(_03301_),
    .X(_03315_));
 sky130_fd_sc_hd__clkbuf_1 _18289_ (.A(_03315_),
    .X(_00347_));
 sky130_fd_sc_hd__nand2_1 _18290_ (.A(_03312_),
    .B(_12198_),
    .Y(_03316_));
 sky130_fd_sc_hd__o211a_1 _18291_ (.A1(_03228_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_1 _18292_ (.A0(_03317_),
    .A1(net2019),
    .S(_03301_),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _18293_ (.A(_03318_),
    .X(_00348_));
 sky130_fd_sc_hd__nand2_1 _18294_ (.A(_03312_),
    .B(_12206_),
    .Y(_03319_));
 sky130_fd_sc_hd__o211a_1 _18295_ (.A1(_03232_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _18296_ (.A0(_03320_),
    .A1(net2088),
    .S(_03301_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _18297_ (.A(_03321_),
    .X(_00349_));
 sky130_fd_sc_hd__nand2_1 _18298_ (.A(_03312_),
    .B(_12214_),
    .Y(_03322_));
 sky130_fd_sc_hd__o211a_1 _18299_ (.A1(_03236_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _18300_ (.A0(_03323_),
    .A1(net2113),
    .S(_03301_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_1 _18301_ (.A(_03324_),
    .X(_00350_));
 sky130_fd_sc_hd__nand2_1 _18302_ (.A(_03312_),
    .B(_12222_),
    .Y(_03325_));
 sky130_fd_sc_hd__o211a_1 _18303_ (.A1(_03240_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_1 _18304_ (.A0(_03326_),
    .A1(net2274),
    .S(_03301_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_1 _18305_ (.A(_03327_),
    .X(_00351_));
 sky130_fd_sc_hd__nand2_1 _18306_ (.A(_03312_),
    .B(_12230_),
    .Y(_03328_));
 sky130_fd_sc_hd__o211a_1 _18307_ (.A1(_03244_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _18308_ (.A0(_03329_),
    .A1(net2101),
    .S(_03301_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _18309_ (.A(_03330_),
    .X(_00352_));
 sky130_fd_sc_hd__nand2_1 _18310_ (.A(_03312_),
    .B(_12238_),
    .Y(_03331_));
 sky130_fd_sc_hd__o211a_1 _18311_ (.A1(_03248_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _18312_ (.A0(_03332_),
    .A1(net2199),
    .S(_03301_),
    .X(_03333_));
 sky130_fd_sc_hd__clkbuf_1 _18313_ (.A(_03333_),
    .X(_00353_));
 sky130_fd_sc_hd__nand2_1 _18314_ (.A(_03312_),
    .B(_12246_),
    .Y(_03334_));
 sky130_fd_sc_hd__o211a_1 _18315_ (.A1(_03252_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _18316_ (.A0(_03335_),
    .A1(net2034),
    .S(_03301_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _18317_ (.A(_03336_),
    .X(_00354_));
 sky130_fd_sc_hd__o211a_1 _18318_ (.A1(_03256_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03313_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_8 _18319_ (.A(_03300_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _18320_ (.A0(_03337_),
    .A1(net2270),
    .S(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__clkbuf_1 _18321_ (.A(_03339_),
    .X(_00355_));
 sky130_fd_sc_hd__o211a_1 _18322_ (.A1(_03261_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03316_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _18323_ (.A0(_03340_),
    .A1(net2920),
    .S(_03338_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_1 _18324_ (.A(_03341_),
    .X(_00356_));
 sky130_fd_sc_hd__o211a_1 _18325_ (.A1(_03264_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03319_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _18326_ (.A0(_03342_),
    .A1(net2356),
    .S(_03338_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _18327_ (.A(_03343_),
    .X(_00357_));
 sky130_fd_sc_hd__o211a_1 _18328_ (.A1(_03267_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03322_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _18329_ (.A0(_03344_),
    .A1(net3500),
    .S(_03338_),
    .X(_03345_));
 sky130_fd_sc_hd__clkbuf_1 _18330_ (.A(_03345_),
    .X(_00358_));
 sky130_fd_sc_hd__o211a_1 _18331_ (.A1(_03270_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03325_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _18332_ (.A0(_03346_),
    .A1(net3015),
    .S(_03338_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_1 _18333_ (.A(_03347_),
    .X(_00359_));
 sky130_fd_sc_hd__o211a_1 _18334_ (.A1(_03273_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03328_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _18335_ (.A0(_03348_),
    .A1(net2560),
    .S(_03338_),
    .X(_03349_));
 sky130_fd_sc_hd__clkbuf_1 _18336_ (.A(_03349_),
    .X(_00360_));
 sky130_fd_sc_hd__o211a_1 _18337_ (.A1(_03276_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03331_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _18338_ (.A0(_03350_),
    .A1(net2318),
    .S(_03338_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_1 _18339_ (.A(_03351_),
    .X(_00361_));
 sky130_fd_sc_hd__o211a_1 _18340_ (.A1(_03279_),
    .A2(_03310_),
    .B1(_03311_),
    .C1(_03334_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _18341_ (.A0(_03352_),
    .A1(net2813),
    .S(_03338_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_1 _18342_ (.A(_03353_),
    .X(_00362_));
 sky130_fd_sc_hd__buf_4 _18343_ (.A(_12180_),
    .X(_03354_));
 sky130_fd_sc_hd__o211a_1 _18344_ (.A1(_12170_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03313_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _18345_ (.A0(_03355_),
    .A1(net2531),
    .S(_03338_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _18346_ (.A(_03356_),
    .X(_00363_));
 sky130_fd_sc_hd__o211a_1 _18347_ (.A1(_12195_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03316_),
    .X(_03357_));
 sky130_fd_sc_hd__mux2_1 _18348_ (.A0(_03357_),
    .A1(net2781),
    .S(_03338_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _18349_ (.A(_03358_),
    .X(_00364_));
 sky130_fd_sc_hd__o211a_1 _18350_ (.A1(_12203_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03319_),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_1 _18351_ (.A0(_03359_),
    .A1(net2612),
    .S(_03338_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_1 _18352_ (.A(_03360_),
    .X(_00365_));
 sky130_fd_sc_hd__o211a_1 _18353_ (.A1(_12211_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03322_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _18354_ (.A0(_03361_),
    .A1(net2620),
    .S(_03338_),
    .X(_03362_));
 sky130_fd_sc_hd__clkbuf_1 _18355_ (.A(_03362_),
    .X(_00366_));
 sky130_fd_sc_hd__o211a_1 _18356_ (.A1(_12219_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03325_),
    .X(_03363_));
 sky130_fd_sc_hd__mux2_1 _18357_ (.A0(_03363_),
    .A1(net3481),
    .S(_03338_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _18358_ (.A(_03364_),
    .X(_00367_));
 sky130_fd_sc_hd__o211a_1 _18359_ (.A1(_12227_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03328_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_1 _18360_ (.A0(_03365_),
    .A1(net2828),
    .S(_03338_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_1 _18361_ (.A(_03366_),
    .X(_00368_));
 sky130_fd_sc_hd__o211a_1 _18362_ (.A1(_12235_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03331_),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _18363_ (.A0(_03367_),
    .A1(net2926),
    .S(_03338_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _18364_ (.A(_03368_),
    .X(_00369_));
 sky130_fd_sc_hd__o211a_1 _18365_ (.A1(_12243_),
    .A2(_03312_),
    .B1(_03354_),
    .C1(_03334_),
    .X(_03369_));
 sky130_fd_sc_hd__mux2_1 _18366_ (.A0(_03369_),
    .A1(net3412),
    .S(_03338_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _18367_ (.A(_03370_),
    .X(_00370_));
 sky130_fd_sc_hd__nor2_2 _18368_ (.A(_12292_),
    .B(_03208_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_4 _18369_ (.A(_03371_),
    .B(_12313_),
    .Y(_03372_));
 sky130_fd_sc_hd__a21bo_1 _18370_ (.A1(_03372_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_8 _18371_ (.A(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _18372_ (.A0(_02810_),
    .A1(net2924),
    .S(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _18373_ (.A(_03375_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _18374_ (.A0(_02823_),
    .A1(net3703),
    .S(_03374_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _18375_ (.A(_03376_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _18376_ (.A0(_02827_),
    .A1(net2965),
    .S(_03374_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _18377_ (.A(_03377_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _18378_ (.A0(_02831_),
    .A1(net3669),
    .S(_03374_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _18379_ (.A(_03378_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _18380_ (.A0(_02835_),
    .A1(net3732),
    .S(_03374_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _18381_ (.A(_03379_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _18382_ (.A0(_02839_),
    .A1(net3266),
    .S(_03374_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_1 _18383_ (.A(_03380_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _18384_ (.A0(_02843_),
    .A1(net3208),
    .S(_03374_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_1 _18385_ (.A(_03381_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _18386_ (.A0(_02847_),
    .A1(net3150),
    .S(_03374_),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_1 _18387_ (.A(_03382_),
    .X(_00378_));
 sky130_fd_sc_hd__buf_4 _18388_ (.A(_03372_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_4 _18389_ (.A(_03372_),
    .X(_03384_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(_03384_),
    .B(_12185_),
    .Y(_03385_));
 sky130_fd_sc_hd__o211a_1 _18391_ (.A1(_03222_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _18392_ (.A0(_03386_),
    .A1(net2524),
    .S(_03374_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_1 _18393_ (.A(_03387_),
    .X(_00379_));
 sky130_fd_sc_hd__nand2_1 _18394_ (.A(_03384_),
    .B(_12198_),
    .Y(_03388_));
 sky130_fd_sc_hd__o211a_1 _18395_ (.A1(_03228_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__mux2_1 _18396_ (.A0(_03389_),
    .A1(net3688),
    .S(_03374_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _18397_ (.A(_03390_),
    .X(_00380_));
 sky130_fd_sc_hd__nand2_1 _18398_ (.A(_03384_),
    .B(_12206_),
    .Y(_03391_));
 sky130_fd_sc_hd__o211a_1 _18399_ (.A1(_03232_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _18400_ (.A0(_03392_),
    .A1(net2862),
    .S(_03374_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _18401_ (.A(_03393_),
    .X(_00381_));
 sky130_fd_sc_hd__nand2_1 _18402_ (.A(_03384_),
    .B(_12214_),
    .Y(_03394_));
 sky130_fd_sc_hd__o211a_1 _18403_ (.A1(_03236_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__mux2_1 _18404_ (.A0(_03395_),
    .A1(net3603),
    .S(_03374_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _18405_ (.A(_03396_),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_1 _18406_ (.A(_03384_),
    .B(_12222_),
    .Y(_03397_));
 sky130_fd_sc_hd__o211a_1 _18407_ (.A1(_03240_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _18408_ (.A0(_03398_),
    .A1(net3652),
    .S(_03374_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _18409_ (.A(_03399_),
    .X(_00383_));
 sky130_fd_sc_hd__nand2_1 _18410_ (.A(_03384_),
    .B(_12230_),
    .Y(_03400_));
 sky130_fd_sc_hd__o211a_1 _18411_ (.A1(_03244_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__mux2_1 _18412_ (.A0(_03401_),
    .A1(net2513),
    .S(_03374_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_1 _18413_ (.A(_03402_),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _18414_ (.A(_03384_),
    .B(_12238_),
    .Y(_03403_));
 sky130_fd_sc_hd__o211a_1 _18415_ (.A1(_03248_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_1 _18416_ (.A0(_03404_),
    .A1(net3367),
    .S(_03374_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _18417_ (.A(_03405_),
    .X(_00385_));
 sky130_fd_sc_hd__nand2_1 _18418_ (.A(_03384_),
    .B(_12246_),
    .Y(_03406_));
 sky130_fd_sc_hd__o211a_1 _18419_ (.A1(_03252_),
    .A2(_03383_),
    .B1(_03354_),
    .C1(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__mux2_1 _18420_ (.A0(_03407_),
    .A1(net2735),
    .S(_03374_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _18421_ (.A(_03408_),
    .X(_00386_));
 sky130_fd_sc_hd__buf_4 _18422_ (.A(_12180_),
    .X(_03409_));
 sky130_fd_sc_hd__o211a_1 _18423_ (.A1(_03256_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03385_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_8 _18424_ (.A(_03373_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _18425_ (.A0(_03410_),
    .A1(net2323),
    .S(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _18426_ (.A(_03412_),
    .X(_00387_));
 sky130_fd_sc_hd__o211a_1 _18427_ (.A1(_03261_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03388_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _18428_ (.A0(_03413_),
    .A1(net2536),
    .S(_03411_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _18429_ (.A(_03414_),
    .X(_00388_));
 sky130_fd_sc_hd__o211a_1 _18430_ (.A1(_03264_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03391_),
    .X(_03415_));
 sky130_fd_sc_hd__mux2_1 _18431_ (.A0(_03415_),
    .A1(net2415),
    .S(_03411_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _18432_ (.A(_03416_),
    .X(_00389_));
 sky130_fd_sc_hd__o211a_1 _18433_ (.A1(_03267_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03394_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _18434_ (.A0(_03417_),
    .A1(net2765),
    .S(_03411_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _18435_ (.A(_03418_),
    .X(_00390_));
 sky130_fd_sc_hd__o211a_1 _18436_ (.A1(_03270_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03397_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _18437_ (.A0(_03419_),
    .A1(net2543),
    .S(_03411_),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _18438_ (.A(_03420_),
    .X(_00391_));
 sky130_fd_sc_hd__o211a_1 _18439_ (.A1(_03273_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03400_),
    .X(_03421_));
 sky130_fd_sc_hd__mux2_1 _18440_ (.A0(_03421_),
    .A1(net2643),
    .S(_03411_),
    .X(_03422_));
 sky130_fd_sc_hd__clkbuf_1 _18441_ (.A(_03422_),
    .X(_00392_));
 sky130_fd_sc_hd__o211a_1 _18442_ (.A1(_03276_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03403_),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _18443_ (.A0(_03423_),
    .A1(net2486),
    .S(_03411_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_1 _18444_ (.A(_03424_),
    .X(_00393_));
 sky130_fd_sc_hd__o211a_1 _18445_ (.A1(_03279_),
    .A2(_03383_),
    .B1(_03409_),
    .C1(_03406_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _18446_ (.A0(_03425_),
    .A1(net2405),
    .S(_03411_),
    .X(_03426_));
 sky130_fd_sc_hd__clkbuf_1 _18447_ (.A(_03426_),
    .X(_00394_));
 sky130_fd_sc_hd__o211a_1 _18448_ (.A1(_12170_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03385_),
    .X(_03427_));
 sky130_fd_sc_hd__mux2_1 _18449_ (.A0(_03427_),
    .A1(net2454),
    .S(_03411_),
    .X(_03428_));
 sky130_fd_sc_hd__clkbuf_1 _18450_ (.A(_03428_),
    .X(_00395_));
 sky130_fd_sc_hd__o211a_1 _18451_ (.A1(_12195_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03388_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _18452_ (.A0(_03429_),
    .A1(net2726),
    .S(_03411_),
    .X(_03430_));
 sky130_fd_sc_hd__clkbuf_1 _18453_ (.A(_03430_),
    .X(_00396_));
 sky130_fd_sc_hd__o211a_1 _18454_ (.A1(_12203_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03391_),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_1 _18455_ (.A0(_03431_),
    .A1(net2909),
    .S(_03411_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _18456_ (.A(_03432_),
    .X(_00397_));
 sky130_fd_sc_hd__o211a_1 _18457_ (.A1(_12211_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03394_),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _18458_ (.A0(_03433_),
    .A1(net2604),
    .S(_03411_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _18459_ (.A(_03434_),
    .X(_00398_));
 sky130_fd_sc_hd__o211a_1 _18460_ (.A1(_12219_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03397_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _18461_ (.A0(_03435_),
    .A1(net2736),
    .S(_03411_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _18462_ (.A(_03436_),
    .X(_00399_));
 sky130_fd_sc_hd__o211a_1 _18463_ (.A1(_12227_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03400_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _18464_ (.A0(_03437_),
    .A1(net3463),
    .S(_03411_),
    .X(_03438_));
 sky130_fd_sc_hd__clkbuf_1 _18465_ (.A(_03438_),
    .X(_00400_));
 sky130_fd_sc_hd__o211a_1 _18466_ (.A1(_12235_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03403_),
    .X(_03439_));
 sky130_fd_sc_hd__mux2_1 _18467_ (.A0(_03439_),
    .A1(net2956),
    .S(_03411_),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_1 _18468_ (.A(_03440_),
    .X(_00401_));
 sky130_fd_sc_hd__o211a_1 _18469_ (.A1(_12243_),
    .A2(_03384_),
    .B1(_03409_),
    .C1(_03406_),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_1 _18470_ (.A0(_03441_),
    .A1(net3476),
    .S(_03411_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_1 _18471_ (.A(_03442_),
    .X(_00402_));
 sky130_fd_sc_hd__nor2_1 _18472_ (.A(_12171_),
    .B(_03208_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2_4 _18473_ (.A(_03443_),
    .B(_12313_),
    .Y(_03444_));
 sky130_fd_sc_hd__a21bo_1 _18474_ (.A1(_03444_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_8 _18475_ (.A(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__mux2_1 _18476_ (.A0(_02810_),
    .A1(net2622),
    .S(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _18477_ (.A(_03447_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _18478_ (.A0(_02823_),
    .A1(net2973),
    .S(_03446_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_1 _18479_ (.A(_03448_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _18480_ (.A0(_02827_),
    .A1(net3170),
    .S(_03446_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_1 _18481_ (.A(_03449_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _18482_ (.A0(_02831_),
    .A1(net2928),
    .S(_03446_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _18483_ (.A(_03450_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _18484_ (.A0(_02835_),
    .A1(net3487),
    .S(_03446_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _18485_ (.A(_03451_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _18486_ (.A0(_02839_),
    .A1(net2477),
    .S(_03446_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_1 _18487_ (.A(_03452_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _18488_ (.A0(_02843_),
    .A1(net2269),
    .S(_03446_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _18489_ (.A(_03453_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _18490_ (.A0(_02847_),
    .A1(net3274),
    .S(_03446_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_1 _18491_ (.A(_03454_),
    .X(_00410_));
 sky130_fd_sc_hd__buf_4 _18492_ (.A(_03444_),
    .X(_03455_));
 sky130_fd_sc_hd__buf_4 _18493_ (.A(_12180_),
    .X(_03456_));
 sky130_fd_sc_hd__buf_4 _18494_ (.A(_03444_),
    .X(_03457_));
 sky130_fd_sc_hd__nand2_1 _18495_ (.A(_03457_),
    .B(_12185_),
    .Y(_03458_));
 sky130_fd_sc_hd__o211a_1 _18496_ (.A1(_03222_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _18497_ (.A0(_03459_),
    .A1(net2796),
    .S(_03446_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _18498_ (.A(_03460_),
    .X(_00411_));
 sky130_fd_sc_hd__nand2_1 _18499_ (.A(_03457_),
    .B(_12198_),
    .Y(_03461_));
 sky130_fd_sc_hd__o211a_1 _18500_ (.A1(_03228_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__mux2_1 _18501_ (.A0(_03462_),
    .A1(net3010),
    .S(_03446_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _18502_ (.A(_03463_),
    .X(_00412_));
 sky130_fd_sc_hd__nand2_1 _18503_ (.A(_03457_),
    .B(_12206_),
    .Y(_03464_));
 sky130_fd_sc_hd__o211a_1 _18504_ (.A1(_03232_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__mux2_1 _18505_ (.A0(_03465_),
    .A1(net2811),
    .S(_03446_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _18506_ (.A(_03466_),
    .X(_00413_));
 sky130_fd_sc_hd__nand2_1 _18507_ (.A(_03457_),
    .B(_12214_),
    .Y(_03467_));
 sky130_fd_sc_hd__o211a_1 _18508_ (.A1(_03236_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_1 _18509_ (.A0(_03468_),
    .A1(net3275),
    .S(_03446_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _18510_ (.A(_03469_),
    .X(_00414_));
 sky130_fd_sc_hd__nand2_1 _18511_ (.A(_03457_),
    .B(_12222_),
    .Y(_03470_));
 sky130_fd_sc_hd__o211a_1 _18512_ (.A1(_03240_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__mux2_1 _18513_ (.A0(_03471_),
    .A1(net2687),
    .S(_03446_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _18514_ (.A(_03472_),
    .X(_00415_));
 sky130_fd_sc_hd__nand2_1 _18515_ (.A(_03457_),
    .B(_12230_),
    .Y(_03473_));
 sky130_fd_sc_hd__o211a_1 _18516_ (.A1(_03244_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _18517_ (.A0(_03474_),
    .A1(net2891),
    .S(_03446_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _18518_ (.A(_03475_),
    .X(_00416_));
 sky130_fd_sc_hd__nand2_1 _18519_ (.A(_03457_),
    .B(_12238_),
    .Y(_03476_));
 sky130_fd_sc_hd__o211a_1 _18520_ (.A1(_03248_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_1 _18521_ (.A0(_03477_),
    .A1(net2453),
    .S(_03446_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _18522_ (.A(_03478_),
    .X(_00417_));
 sky130_fd_sc_hd__nand2_1 _18523_ (.A(_03457_),
    .B(_12246_),
    .Y(_03479_));
 sky130_fd_sc_hd__o211a_1 _18524_ (.A1(_03252_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _18525_ (.A0(_03480_),
    .A1(net2818),
    .S(_03446_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_1 _18526_ (.A(_03481_),
    .X(_00418_));
 sky130_fd_sc_hd__o211a_1 _18527_ (.A1(_03256_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03458_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_8 _18528_ (.A(_03445_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _18529_ (.A0(_03482_),
    .A1(net2901),
    .S(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _18530_ (.A(_03484_),
    .X(_00419_));
 sky130_fd_sc_hd__o211a_1 _18531_ (.A1(_03261_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03461_),
    .X(_03485_));
 sky130_fd_sc_hd__mux2_1 _18532_ (.A0(_03485_),
    .A1(net2313),
    .S(_03483_),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_1 _18533_ (.A(_03486_),
    .X(_00420_));
 sky130_fd_sc_hd__o211a_1 _18534_ (.A1(_03264_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03464_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _18535_ (.A0(_03487_),
    .A1(net3194),
    .S(_03483_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _18536_ (.A(_03488_),
    .X(_00421_));
 sky130_fd_sc_hd__o211a_1 _18537_ (.A1(_03267_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03467_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _18538_ (.A0(_03489_),
    .A1(net2708),
    .S(_03483_),
    .X(_03490_));
 sky130_fd_sc_hd__clkbuf_1 _18539_ (.A(_03490_),
    .X(_00422_));
 sky130_fd_sc_hd__o211a_1 _18540_ (.A1(_03270_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03470_),
    .X(_03491_));
 sky130_fd_sc_hd__mux2_1 _18541_ (.A0(_03491_),
    .A1(net2880),
    .S(_03483_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _18542_ (.A(_03492_),
    .X(_00423_));
 sky130_fd_sc_hd__o211a_1 _18543_ (.A1(_03273_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03473_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_1 _18544_ (.A0(_03493_),
    .A1(net2911),
    .S(_03483_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _18545_ (.A(_03494_),
    .X(_00424_));
 sky130_fd_sc_hd__o211a_1 _18546_ (.A1(_03276_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03476_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _18547_ (.A0(_03495_),
    .A1(net2830),
    .S(_03483_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_1 _18548_ (.A(_03496_),
    .X(_00425_));
 sky130_fd_sc_hd__o211a_1 _18549_ (.A1(_03279_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03479_),
    .X(_03497_));
 sky130_fd_sc_hd__mux2_1 _18550_ (.A0(_03497_),
    .A1(net3523),
    .S(_03483_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_1 _18551_ (.A(_03498_),
    .X(_00426_));
 sky130_fd_sc_hd__buf_4 _18552_ (.A(_12180_),
    .X(_03499_));
 sky130_fd_sc_hd__o211a_1 _18553_ (.A1(_12170_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03458_),
    .X(_03500_));
 sky130_fd_sc_hd__mux2_1 _18554_ (.A0(_03500_),
    .A1(net3851),
    .S(_03483_),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_1 _18555_ (.A(_03501_),
    .X(_00427_));
 sky130_fd_sc_hd__o211a_1 _18556_ (.A1(_12195_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03461_),
    .X(_03502_));
 sky130_fd_sc_hd__mux2_1 _18557_ (.A0(_03502_),
    .A1(net3825),
    .S(_03483_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_1 _18558_ (.A(_03503_),
    .X(_00428_));
 sky130_fd_sc_hd__o211a_1 _18559_ (.A1(_12203_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03464_),
    .X(_03504_));
 sky130_fd_sc_hd__mux2_1 _18560_ (.A0(_03504_),
    .A1(net3833),
    .S(_03483_),
    .X(_03505_));
 sky130_fd_sc_hd__clkbuf_1 _18561_ (.A(_03505_),
    .X(_00429_));
 sky130_fd_sc_hd__o211a_1 _18562_ (.A1(_12211_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03467_),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_1 _18563_ (.A0(_03506_),
    .A1(net3845),
    .S(_03483_),
    .X(_03507_));
 sky130_fd_sc_hd__clkbuf_1 _18564_ (.A(_03507_),
    .X(_00430_));
 sky130_fd_sc_hd__o211a_1 _18565_ (.A1(_12219_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03470_),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_1 _18566_ (.A0(_03508_),
    .A1(net3544),
    .S(_03483_),
    .X(_03509_));
 sky130_fd_sc_hd__clkbuf_1 _18567_ (.A(_03509_),
    .X(_00431_));
 sky130_fd_sc_hd__o211a_1 _18568_ (.A1(_12227_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03473_),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_1 _18569_ (.A0(_03510_),
    .A1(net3849),
    .S(_03483_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _18570_ (.A(_03511_),
    .X(_00432_));
 sky130_fd_sc_hd__o211a_1 _18571_ (.A1(_12235_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03476_),
    .X(_03512_));
 sky130_fd_sc_hd__mux2_1 _18572_ (.A0(_03512_),
    .A1(net3808),
    .S(_03483_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_1 _18573_ (.A(_03513_),
    .X(_00433_));
 sky130_fd_sc_hd__o211a_1 _18574_ (.A1(_12243_),
    .A2(_03457_),
    .B1(_03499_),
    .C1(_03479_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _18575_ (.A0(_03514_),
    .A1(net3899),
    .S(_03483_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _18576_ (.A(_03515_),
    .X(_00434_));
 sky130_fd_sc_hd__nor2_2 _18577_ (.A(\line_cache_idx[4] ),
    .B(_09092_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_2 _18578_ (.A(_03516_),
    .B(_12174_),
    .Y(_03517_));
 sky130_fd_sc_hd__or2_1 _18579_ (.A(_02812_),
    .B(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__inv_2 _18580_ (.A(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__nand2_4 _18581_ (.A(_03519_),
    .B(_12313_),
    .Y(_03520_));
 sky130_fd_sc_hd__a21bo_1 _18582_ (.A1(_03520_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03521_));
 sky130_fd_sc_hd__buf_6 _18583_ (.A(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_1 _18584_ (.A0(_02810_),
    .A1(net3453),
    .S(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _18585_ (.A(_03523_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _18586_ (.A0(_02823_),
    .A1(net2883),
    .S(_03522_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _18587_ (.A(_03524_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _18588_ (.A0(_02827_),
    .A1(net2338),
    .S(_03522_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _18589_ (.A(_03525_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _18590_ (.A0(_02831_),
    .A1(net3018),
    .S(_03522_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _18591_ (.A(_03526_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _18592_ (.A0(_02835_),
    .A1(net2345),
    .S(_03522_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _18593_ (.A(_03527_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _18594_ (.A0(_02839_),
    .A1(net3277),
    .S(_03522_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _18595_ (.A(_03528_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _18596_ (.A0(_02843_),
    .A1(net3108),
    .S(_03522_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _18597_ (.A(_03529_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _18598_ (.A0(_02847_),
    .A1(net3068),
    .S(_03522_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _18599_ (.A(_03530_),
    .X(_00442_));
 sky130_fd_sc_hd__buf_4 _18600_ (.A(_03520_),
    .X(_03531_));
 sky130_fd_sc_hd__buf_4 _18601_ (.A(_03520_),
    .X(_03532_));
 sky130_fd_sc_hd__nand2_1 _18602_ (.A(_03532_),
    .B(_12185_),
    .Y(_03533_));
 sky130_fd_sc_hd__o211a_1 _18603_ (.A1(_03222_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _18604_ (.A0(_03534_),
    .A1(net2359),
    .S(_03522_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _18605_ (.A(_03535_),
    .X(_00443_));
 sky130_fd_sc_hd__nand2_1 _18606_ (.A(_03532_),
    .B(_12198_),
    .Y(_03536_));
 sky130_fd_sc_hd__o211a_1 _18607_ (.A1(_03228_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_1 _18608_ (.A0(_03537_),
    .A1(net2654),
    .S(_03522_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _18609_ (.A(_03538_),
    .X(_00444_));
 sky130_fd_sc_hd__nand2_1 _18610_ (.A(_03532_),
    .B(_12206_),
    .Y(_03539_));
 sky130_fd_sc_hd__o211a_1 _18611_ (.A1(_03232_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_1 _18612_ (.A0(_03540_),
    .A1(net2570),
    .S(_03522_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _18613_ (.A(_03541_),
    .X(_00445_));
 sky130_fd_sc_hd__nand2_1 _18614_ (.A(_03532_),
    .B(_12214_),
    .Y(_03542_));
 sky130_fd_sc_hd__o211a_1 _18615_ (.A1(_03236_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _18616_ (.A0(_03543_),
    .A1(net2919),
    .S(_03522_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _18617_ (.A(_03544_),
    .X(_00446_));
 sky130_fd_sc_hd__nand2_1 _18618_ (.A(_03532_),
    .B(_12222_),
    .Y(_03545_));
 sky130_fd_sc_hd__o211a_1 _18619_ (.A1(_03240_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _18620_ (.A0(_03546_),
    .A1(net3441),
    .S(_03522_),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _18621_ (.A(_03547_),
    .X(_00447_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(_03532_),
    .B(_12230_),
    .Y(_03548_));
 sky130_fd_sc_hd__o211a_1 _18623_ (.A1(_03244_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _18624_ (.A0(_03549_),
    .A1(net3041),
    .S(_03522_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _18625_ (.A(_03550_),
    .X(_00448_));
 sky130_fd_sc_hd__nand2_1 _18626_ (.A(_03532_),
    .B(_12238_),
    .Y(_03551_));
 sky130_fd_sc_hd__o211a_1 _18627_ (.A1(_03248_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _18628_ (.A0(_03552_),
    .A1(net2800),
    .S(_03522_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _18629_ (.A(_03553_),
    .X(_00449_));
 sky130_fd_sc_hd__nand2_1 _18630_ (.A(_03532_),
    .B(_12246_),
    .Y(_03554_));
 sky130_fd_sc_hd__o211a_1 _18631_ (.A1(_03252_),
    .A2(_03531_),
    .B1(_03499_),
    .C1(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_1 _18632_ (.A0(_03555_),
    .A1(net2848),
    .S(_03522_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _18633_ (.A(_03556_),
    .X(_00450_));
 sky130_fd_sc_hd__buf_4 _18634_ (.A(_12180_),
    .X(_03557_));
 sky130_fd_sc_hd__o211a_1 _18635_ (.A1(_03256_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03533_),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_8 _18636_ (.A(_03521_),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_1 _18637_ (.A0(_03558_),
    .A1(net2672),
    .S(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _18638_ (.A(_03560_),
    .X(_00451_));
 sky130_fd_sc_hd__o211a_1 _18639_ (.A1(_03261_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03536_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _18640_ (.A0(_03561_),
    .A1(net3475),
    .S(_03559_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _18641_ (.A(_03562_),
    .X(_00452_));
 sky130_fd_sc_hd__o211a_1 _18642_ (.A1(_03264_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03539_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _18643_ (.A0(_03563_),
    .A1(net3088),
    .S(_03559_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _18644_ (.A(_03564_),
    .X(_00453_));
 sky130_fd_sc_hd__o211a_1 _18645_ (.A1(_03267_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03542_),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_1 _18646_ (.A0(_03565_),
    .A1(net3202),
    .S(_03559_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _18647_ (.A(_03566_),
    .X(_00454_));
 sky130_fd_sc_hd__o211a_1 _18648_ (.A1(_03270_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03545_),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_1 _18649_ (.A0(_03567_),
    .A1(net3192),
    .S(_03559_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_1 _18650_ (.A(_03568_),
    .X(_00455_));
 sky130_fd_sc_hd__o211a_1 _18651_ (.A1(_03273_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03548_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _18652_ (.A0(_03569_),
    .A1(net2343),
    .S(_03559_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _18653_ (.A(_03570_),
    .X(_00456_));
 sky130_fd_sc_hd__o211a_1 _18654_ (.A1(_03276_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03551_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _18655_ (.A0(_03571_),
    .A1(net3285),
    .S(_03559_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _18656_ (.A(_03572_),
    .X(_00457_));
 sky130_fd_sc_hd__o211a_1 _18657_ (.A1(_03279_),
    .A2(_03531_),
    .B1(_03557_),
    .C1(_03554_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _18658_ (.A0(_03573_),
    .A1(net3284),
    .S(_03559_),
    .X(_03574_));
 sky130_fd_sc_hd__clkbuf_1 _18659_ (.A(_03574_),
    .X(_00458_));
 sky130_fd_sc_hd__o211a_1 _18660_ (.A1(_12170_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03533_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _18661_ (.A0(_03575_),
    .A1(net3409),
    .S(_03559_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _18662_ (.A(_03576_),
    .X(_00459_));
 sky130_fd_sc_hd__o211a_1 _18663_ (.A1(_12195_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03536_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _18664_ (.A0(_03577_),
    .A1(net2601),
    .S(_03559_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_1 _18665_ (.A(_03578_),
    .X(_00460_));
 sky130_fd_sc_hd__o211a_1 _18666_ (.A1(_12203_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03539_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_1 _18667_ (.A0(_03579_),
    .A1(net2793),
    .S(_03559_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_1 _18668_ (.A(_03580_),
    .X(_00461_));
 sky130_fd_sc_hd__o211a_1 _18669_ (.A1(_12211_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03542_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _18670_ (.A0(_03581_),
    .A1(net2812),
    .S(_03559_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _18671_ (.A(_03582_),
    .X(_00462_));
 sky130_fd_sc_hd__o211a_1 _18672_ (.A1(_12219_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03545_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _18673_ (.A0(_03583_),
    .A1(net2723),
    .S(_03559_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _18674_ (.A(_03584_),
    .X(_00463_));
 sky130_fd_sc_hd__o211a_1 _18675_ (.A1(_12227_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03548_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _18676_ (.A0(_03585_),
    .A1(net3082),
    .S(_03559_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _18677_ (.A(_03586_),
    .X(_00464_));
 sky130_fd_sc_hd__o211a_1 _18678_ (.A1(_12235_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03551_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _18679_ (.A0(_03587_),
    .A1(net3203),
    .S(_03559_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _18680_ (.A(_03588_),
    .X(_00465_));
 sky130_fd_sc_hd__o211a_1 _18681_ (.A1(_12243_),
    .A2(_03532_),
    .B1(_03557_),
    .C1(_03554_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _18682_ (.A0(_03589_),
    .A1(net2771),
    .S(_03559_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _18683_ (.A(_03590_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_2 _18684_ (.A(_12293_),
    .B(_03517_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand2_4 _18685_ (.A(_03591_),
    .B(_12313_),
    .Y(_03592_));
 sky130_fd_sc_hd__a21bo_1 _18686_ (.A1(_03592_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03593_));
 sky130_fd_sc_hd__buf_6 _18687_ (.A(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__mux2_1 _18688_ (.A0(_02810_),
    .A1(net2860),
    .S(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _18689_ (.A(_03595_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _18690_ (.A0(_02823_),
    .A1(net2468),
    .S(_03594_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _18691_ (.A(_03596_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _18692_ (.A0(_02827_),
    .A1(net2799),
    .S(_03594_),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _18693_ (.A(_03597_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _18694_ (.A0(_02831_),
    .A1(net3187),
    .S(_03594_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _18695_ (.A(_03598_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _18696_ (.A0(_02835_),
    .A1(net2929),
    .S(_03594_),
    .X(_03599_));
 sky130_fd_sc_hd__clkbuf_1 _18697_ (.A(_03599_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _18698_ (.A0(_02839_),
    .A1(net3126),
    .S(_03594_),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _18699_ (.A(_03600_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _18700_ (.A0(_02843_),
    .A1(net3322),
    .S(_03594_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _18701_ (.A(_03601_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _18702_ (.A0(_02847_),
    .A1(net3280),
    .S(_03594_),
    .X(_03602_));
 sky130_fd_sc_hd__clkbuf_1 _18703_ (.A(_03602_),
    .X(_00474_));
 sky130_fd_sc_hd__buf_4 _18704_ (.A(_03592_),
    .X(_03603_));
 sky130_fd_sc_hd__buf_4 _18705_ (.A(_12180_),
    .X(_03604_));
 sky130_fd_sc_hd__buf_4 _18706_ (.A(_03592_),
    .X(_03605_));
 sky130_fd_sc_hd__nand2_1 _18707_ (.A(_03605_),
    .B(_12185_),
    .Y(_03606_));
 sky130_fd_sc_hd__o211a_1 _18708_ (.A1(_03222_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _18709_ (.A0(_03607_),
    .A1(net2293),
    .S(_03594_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _18710_ (.A(_03608_),
    .X(_00475_));
 sky130_fd_sc_hd__nand2_1 _18711_ (.A(_03605_),
    .B(_12198_),
    .Y(_03609_));
 sky130_fd_sc_hd__o211a_1 _18712_ (.A1(_03228_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _18713_ (.A0(_03610_),
    .A1(net2208),
    .S(_03594_),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _18714_ (.A(_03611_),
    .X(_00476_));
 sky130_fd_sc_hd__nand2_1 _18715_ (.A(_03605_),
    .B(_12206_),
    .Y(_03612_));
 sky130_fd_sc_hd__o211a_1 _18716_ (.A1(_03232_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _18717_ (.A0(_03613_),
    .A1(net2243),
    .S(_03594_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_1 _18718_ (.A(_03614_),
    .X(_00477_));
 sky130_fd_sc_hd__nand2_1 _18719_ (.A(_03605_),
    .B(_12214_),
    .Y(_03615_));
 sky130_fd_sc_hd__o211a_1 _18720_ (.A1(_03236_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _18721_ (.A0(_03616_),
    .A1(net2825),
    .S(_03594_),
    .X(_03617_));
 sky130_fd_sc_hd__clkbuf_1 _18722_ (.A(_03617_),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_1 _18723_ (.A(_03605_),
    .B(_12222_),
    .Y(_03618_));
 sky130_fd_sc_hd__o211a_1 _18724_ (.A1(_03240_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_1 _18725_ (.A0(_03619_),
    .A1(net2462),
    .S(_03594_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _18726_ (.A(_03620_),
    .X(_00479_));
 sky130_fd_sc_hd__nand2_1 _18727_ (.A(_03605_),
    .B(_12230_),
    .Y(_03621_));
 sky130_fd_sc_hd__o211a_1 _18728_ (.A1(_03244_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _18729_ (.A0(_03622_),
    .A1(net2499),
    .S(_03594_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _18730_ (.A(_03623_),
    .X(_00480_));
 sky130_fd_sc_hd__nand2_1 _18731_ (.A(_03605_),
    .B(_12238_),
    .Y(_03624_));
 sky130_fd_sc_hd__o211a_1 _18732_ (.A1(_03248_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _18733_ (.A0(_03625_),
    .A1(net2265),
    .S(_03594_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _18734_ (.A(_03626_),
    .X(_00481_));
 sky130_fd_sc_hd__nand2_1 _18735_ (.A(_03605_),
    .B(_12246_),
    .Y(_03627_));
 sky130_fd_sc_hd__o211a_1 _18736_ (.A1(_03252_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _18737_ (.A0(_03628_),
    .A1(net2824),
    .S(_03594_),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _18738_ (.A(_03629_),
    .X(_00482_));
 sky130_fd_sc_hd__o211a_1 _18739_ (.A1(_03256_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03606_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_8 _18740_ (.A(_03593_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _18741_ (.A0(_03630_),
    .A1(net2239),
    .S(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _18742_ (.A(_03632_),
    .X(_00483_));
 sky130_fd_sc_hd__o211a_1 _18743_ (.A1(_03261_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03609_),
    .X(_03633_));
 sky130_fd_sc_hd__mux2_1 _18744_ (.A0(_03633_),
    .A1(net2440),
    .S(_03631_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_1 _18745_ (.A(_03634_),
    .X(_00484_));
 sky130_fd_sc_hd__o211a_1 _18746_ (.A1(_03264_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03612_),
    .X(_03635_));
 sky130_fd_sc_hd__mux2_1 _18747_ (.A0(_03635_),
    .A1(net2185),
    .S(_03631_),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_1 _18748_ (.A(_03636_),
    .X(_00485_));
 sky130_fd_sc_hd__o211a_1 _18749_ (.A1(_03267_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03615_),
    .X(_03637_));
 sky130_fd_sc_hd__mux2_1 _18750_ (.A0(_03637_),
    .A1(net2768),
    .S(_03631_),
    .X(_03638_));
 sky130_fd_sc_hd__clkbuf_1 _18751_ (.A(_03638_),
    .X(_00486_));
 sky130_fd_sc_hd__o211a_1 _18752_ (.A1(_03270_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03618_),
    .X(_03639_));
 sky130_fd_sc_hd__mux2_1 _18753_ (.A0(_03639_),
    .A1(net2283),
    .S(_03631_),
    .X(_03640_));
 sky130_fd_sc_hd__clkbuf_1 _18754_ (.A(_03640_),
    .X(_00487_));
 sky130_fd_sc_hd__o211a_1 _18755_ (.A1(_03273_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03621_),
    .X(_03641_));
 sky130_fd_sc_hd__mux2_1 _18756_ (.A0(_03641_),
    .A1(net2671),
    .S(_03631_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_1 _18757_ (.A(_03642_),
    .X(_00488_));
 sky130_fd_sc_hd__o211a_1 _18758_ (.A1(_03276_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03624_),
    .X(_03643_));
 sky130_fd_sc_hd__mux2_1 _18759_ (.A0(_03643_),
    .A1(net3407),
    .S(_03631_),
    .X(_03644_));
 sky130_fd_sc_hd__clkbuf_1 _18760_ (.A(_03644_),
    .X(_00489_));
 sky130_fd_sc_hd__o211a_1 _18761_ (.A1(_03279_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03627_),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_1 _18762_ (.A0(_03645_),
    .A1(net2806),
    .S(_03631_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_1 _18763_ (.A(_03646_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_4 _18764_ (.A(_12180_),
    .X(_03647_));
 sky130_fd_sc_hd__o211a_1 _18765_ (.A1(_12170_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03606_),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _18766_ (.A0(_03648_),
    .A1(net3680),
    .S(_03631_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _18767_ (.A(_03649_),
    .X(_00491_));
 sky130_fd_sc_hd__o211a_1 _18768_ (.A1(_12195_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03609_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _18769_ (.A0(_03650_),
    .A1(net3565),
    .S(_03631_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _18770_ (.A(_03651_),
    .X(_00492_));
 sky130_fd_sc_hd__o211a_1 _18771_ (.A1(_12203_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03612_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _18772_ (.A0(_03652_),
    .A1(net2910),
    .S(_03631_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_1 _18773_ (.A(_03653_),
    .X(_00493_));
 sky130_fd_sc_hd__o211a_1 _18774_ (.A1(_12211_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03615_),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _18775_ (.A0(_03654_),
    .A1(net3668),
    .S(_03631_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_1 _18776_ (.A(_03655_),
    .X(_00494_));
 sky130_fd_sc_hd__o211a_1 _18777_ (.A1(_12219_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03618_),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _18778_ (.A0(_03656_),
    .A1(net3712),
    .S(_03631_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _18779_ (.A(_03657_),
    .X(_00495_));
 sky130_fd_sc_hd__o211a_1 _18780_ (.A1(_12227_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03621_),
    .X(_03658_));
 sky130_fd_sc_hd__mux2_1 _18781_ (.A0(_03658_),
    .A1(net3875),
    .S(_03631_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_1 _18782_ (.A(_03659_),
    .X(_00496_));
 sky130_fd_sc_hd__o211a_1 _18783_ (.A1(_12235_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03624_),
    .X(_03660_));
 sky130_fd_sc_hd__mux2_1 _18784_ (.A0(_03660_),
    .A1(net3878),
    .S(_03631_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_1 _18785_ (.A(_03661_),
    .X(_00497_));
 sky130_fd_sc_hd__o211a_1 _18786_ (.A1(_12243_),
    .A2(_03605_),
    .B1(_03647_),
    .C1(_03627_),
    .X(_03662_));
 sky130_fd_sc_hd__mux2_1 _18787_ (.A0(_03662_),
    .A1(net3696),
    .S(_03631_),
    .X(_03663_));
 sky130_fd_sc_hd__clkbuf_1 _18788_ (.A(_03663_),
    .X(_00498_));
 sky130_fd_sc_hd__nor2_1 _18789_ (.A(_12292_),
    .B(_03517_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand2_4 _18790_ (.A(_03664_),
    .B(_12313_),
    .Y(_03665_));
 sky130_fd_sc_hd__a21bo_1 _18791_ (.A1(_03665_),
    .A2(_09110_),
    .B1_N(_12190_),
    .X(_03666_));
 sky130_fd_sc_hd__buf_6 _18792_ (.A(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _18793_ (.A0(_02810_),
    .A1(net3681),
    .S(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _18794_ (.A(_03668_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _18795_ (.A0(_02823_),
    .A1(net3705),
    .S(_03667_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _18796_ (.A(_03669_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _18797_ (.A0(_02827_),
    .A1(net2507),
    .S(_03667_),
    .X(_03670_));
 sky130_fd_sc_hd__clkbuf_1 _18798_ (.A(_03670_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _18799_ (.A0(_02831_),
    .A1(net3694),
    .S(_03667_),
    .X(_03671_));
 sky130_fd_sc_hd__clkbuf_1 _18800_ (.A(_03671_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _18801_ (.A0(_02835_),
    .A1(net3741),
    .S(_03667_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _18802_ (.A(_03672_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _18803_ (.A0(_02839_),
    .A1(net3912),
    .S(_03667_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _18804_ (.A(_03673_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _18805_ (.A0(_02843_),
    .A1(net3882),
    .S(_03667_),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_1 _18806_ (.A(_03674_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _18807_ (.A0(_02847_),
    .A1(net3767),
    .S(_03667_),
    .X(_03675_));
 sky130_fd_sc_hd__clkbuf_1 _18808_ (.A(_03675_),
    .X(_00506_));
 sky130_fd_sc_hd__buf_4 _18809_ (.A(_03665_),
    .X(_03676_));
 sky130_fd_sc_hd__buf_4 _18810_ (.A(_03665_),
    .X(_03677_));
 sky130_fd_sc_hd__nand2_1 _18811_ (.A(_03677_),
    .B(_12185_),
    .Y(_03678_));
 sky130_fd_sc_hd__o211a_1 _18812_ (.A1(_03222_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _18813_ (.A0(_03679_),
    .A1(net2168),
    .S(_03667_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _18814_ (.A(_03680_),
    .X(_00507_));
 sky130_fd_sc_hd__nand2_1 _18815_ (.A(_03677_),
    .B(_12198_),
    .Y(_03681_));
 sky130_fd_sc_hd__o211a_1 _18816_ (.A1(_03228_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _18817_ (.A0(_03682_),
    .A1(net2358),
    .S(_03667_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _18818_ (.A(_03683_),
    .X(_00508_));
 sky130_fd_sc_hd__nand2_1 _18819_ (.A(_03677_),
    .B(_12206_),
    .Y(_03684_));
 sky130_fd_sc_hd__o211a_1 _18820_ (.A1(_03232_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _18821_ (.A0(_03685_),
    .A1(net2451),
    .S(_03667_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _18822_ (.A(_03686_),
    .X(_00509_));
 sky130_fd_sc_hd__nand2_1 _18823_ (.A(_03677_),
    .B(_12214_),
    .Y(_03687_));
 sky130_fd_sc_hd__o211a_1 _18824_ (.A1(_03236_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _18825_ (.A0(_03688_),
    .A1(net3014),
    .S(_03667_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _18826_ (.A(_03689_),
    .X(_00510_));
 sky130_fd_sc_hd__nand2_1 _18827_ (.A(_03677_),
    .B(_12222_),
    .Y(_03690_));
 sky130_fd_sc_hd__o211a_1 _18828_ (.A1(_03240_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _18829_ (.A0(_03691_),
    .A1(net2679),
    .S(_03667_),
    .X(_03692_));
 sky130_fd_sc_hd__clkbuf_1 _18830_ (.A(_03692_),
    .X(_00511_));
 sky130_fd_sc_hd__nand2_1 _18831_ (.A(_03677_),
    .B(_12230_),
    .Y(_03693_));
 sky130_fd_sc_hd__o211a_1 _18832_ (.A1(_03244_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _18833_ (.A0(_03694_),
    .A1(net3241),
    .S(_03667_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _18834_ (.A(_03695_),
    .X(_00512_));
 sky130_fd_sc_hd__nand2_1 _18835_ (.A(_03677_),
    .B(_12238_),
    .Y(_03696_));
 sky130_fd_sc_hd__o211a_1 _18836_ (.A1(_03248_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__mux2_1 _18837_ (.A0(_03697_),
    .A1(net2377),
    .S(_03667_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _18838_ (.A(_03698_),
    .X(_00513_));
 sky130_fd_sc_hd__nand2_1 _18839_ (.A(_03677_),
    .B(_12246_),
    .Y(_03699_));
 sky130_fd_sc_hd__o211a_1 _18840_ (.A1(_03252_),
    .A2(_03676_),
    .B1(_03647_),
    .C1(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_1 _18841_ (.A0(_03700_),
    .A1(net2371),
    .S(_03667_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_1 _18842_ (.A(_03701_),
    .X(_00514_));
 sky130_fd_sc_hd__buf_8 _18843_ (.A(_09125_),
    .X(_03702_));
 sky130_fd_sc_hd__buf_4 _18844_ (.A(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__o211a_1 _18845_ (.A1(_03256_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03678_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_8 _18846_ (.A(_03666_),
    .X(_03705_));
 sky130_fd_sc_hd__mux2_1 _18847_ (.A0(_03704_),
    .A1(net2130),
    .S(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_1 _18848_ (.A(_03706_),
    .X(_00515_));
 sky130_fd_sc_hd__o211a_1 _18849_ (.A1(_03261_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03681_),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _18850_ (.A0(_03707_),
    .A1(net2923),
    .S(_03705_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_1 _18851_ (.A(_03708_),
    .X(_00516_));
 sky130_fd_sc_hd__o211a_1 _18852_ (.A1(_03264_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03684_),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_1 _18853_ (.A0(_03709_),
    .A1(net2175),
    .S(_03705_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _18854_ (.A(_03710_),
    .X(_00517_));
 sky130_fd_sc_hd__o211a_1 _18855_ (.A1(_03267_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03687_),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _18856_ (.A0(_03711_),
    .A1(net2223),
    .S(_03705_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_1 _18857_ (.A(_03712_),
    .X(_00518_));
 sky130_fd_sc_hd__o211a_1 _18858_ (.A1(_03270_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03690_),
    .X(_03713_));
 sky130_fd_sc_hd__mux2_1 _18859_ (.A0(_03713_),
    .A1(net2596),
    .S(_03705_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_1 _18860_ (.A(_03714_),
    .X(_00519_));
 sky130_fd_sc_hd__o211a_1 _18861_ (.A1(_03273_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03693_),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_1 _18862_ (.A0(_03715_),
    .A1(net2583),
    .S(_03705_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_1 _18863_ (.A(_03716_),
    .X(_00520_));
 sky130_fd_sc_hd__o211a_1 _18864_ (.A1(_03276_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03696_),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _18865_ (.A0(_03717_),
    .A1(net2339),
    .S(_03705_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_1 _18866_ (.A(_03718_),
    .X(_00521_));
 sky130_fd_sc_hd__o211a_1 _18867_ (.A1(_03279_),
    .A2(_03676_),
    .B1(_03703_),
    .C1(_03699_),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _18868_ (.A0(_03719_),
    .A1(net3129),
    .S(_03705_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _18869_ (.A(_03720_),
    .X(_00522_));
 sky130_fd_sc_hd__o211a_1 _18870_ (.A1(_12170_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03678_),
    .X(_03721_));
 sky130_fd_sc_hd__mux2_1 _18871_ (.A0(_03721_),
    .A1(net3742),
    .S(_03705_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_1 _18872_ (.A(_03722_),
    .X(_00523_));
 sky130_fd_sc_hd__o211a_1 _18873_ (.A1(_12195_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03681_),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_1 _18874_ (.A0(_03723_),
    .A1(net3772),
    .S(_03705_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _18875_ (.A(_03724_),
    .X(_00524_));
 sky130_fd_sc_hd__o211a_1 _18876_ (.A1(_12203_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03684_),
    .X(_03725_));
 sky130_fd_sc_hd__mux2_1 _18877_ (.A0(_03725_),
    .A1(net3892),
    .S(_03705_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_1 _18878_ (.A(_03726_),
    .X(_00525_));
 sky130_fd_sc_hd__o211a_1 _18879_ (.A1(_12211_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03687_),
    .X(_03727_));
 sky130_fd_sc_hd__mux2_1 _18880_ (.A0(_03727_),
    .A1(net3752),
    .S(_03705_),
    .X(_03728_));
 sky130_fd_sc_hd__clkbuf_1 _18881_ (.A(_03728_),
    .X(_00526_));
 sky130_fd_sc_hd__o211a_1 _18882_ (.A1(_12219_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03690_),
    .X(_03729_));
 sky130_fd_sc_hd__mux2_1 _18883_ (.A0(_03729_),
    .A1(net3683),
    .S(_03705_),
    .X(_03730_));
 sky130_fd_sc_hd__clkbuf_1 _18884_ (.A(_03730_),
    .X(_00527_));
 sky130_fd_sc_hd__o211a_1 _18885_ (.A1(_12227_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03693_),
    .X(_03731_));
 sky130_fd_sc_hd__mux2_1 _18886_ (.A0(_03731_),
    .A1(net3676),
    .S(_03705_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_1 _18887_ (.A(_03732_),
    .X(_00528_));
 sky130_fd_sc_hd__o211a_1 _18888_ (.A1(_12235_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03696_),
    .X(_03733_));
 sky130_fd_sc_hd__mux2_1 _18889_ (.A0(_03733_),
    .A1(net3728),
    .S(_03705_),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _18890_ (.A(_03734_),
    .X(_00529_));
 sky130_fd_sc_hd__o211a_1 _18891_ (.A1(_12243_),
    .A2(_03677_),
    .B1(_03703_),
    .C1(_03699_),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_1 _18892_ (.A0(_03735_),
    .A1(net3736),
    .S(_03705_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _18893_ (.A(_03736_),
    .X(_00530_));
 sky130_fd_sc_hd__nor2_1 _18894_ (.A(_12171_),
    .B(_03517_),
    .Y(_03737_));
 sky130_fd_sc_hd__nand2_2 _18895_ (.A(_03737_),
    .B(_12313_),
    .Y(_03738_));
 sky130_fd_sc_hd__buf_12 _18896_ (.A(_12189_),
    .X(_03739_));
 sky130_fd_sc_hd__a21bo_1 _18897_ (.A1(_03738_),
    .A2(_09110_),
    .B1_N(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__buf_6 _18898_ (.A(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _18899_ (.A0(_02810_),
    .A1(net3636),
    .S(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _18900_ (.A(_03742_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _18901_ (.A0(_02823_),
    .A1(net3782),
    .S(_03741_),
    .X(_03743_));
 sky130_fd_sc_hd__clkbuf_1 _18902_ (.A(_03743_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _18903_ (.A0(_02827_),
    .A1(net3871),
    .S(_03741_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _18904_ (.A(_03744_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _18905_ (.A0(_02831_),
    .A1(net3753),
    .S(_03741_),
    .X(_03745_));
 sky130_fd_sc_hd__clkbuf_1 _18906_ (.A(_03745_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _18907_ (.A0(_02835_),
    .A1(net3524),
    .S(_03741_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _18908_ (.A(_03746_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _18909_ (.A0(_02839_),
    .A1(net3550),
    .S(_03741_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _18910_ (.A(_03747_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _18911_ (.A0(_02843_),
    .A1(net3658),
    .S(_03741_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _18912_ (.A(_03748_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _18913_ (.A0(_02847_),
    .A1(net3617),
    .S(_03741_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _18914_ (.A(_03749_),
    .X(_00538_));
 sky130_fd_sc_hd__buf_4 _18915_ (.A(_03738_),
    .X(_03750_));
 sky130_fd_sc_hd__buf_4 _18916_ (.A(_03702_),
    .X(_03751_));
 sky130_fd_sc_hd__buf_4 _18917_ (.A(_03738_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _18918_ (.A(_03752_),
    .B(_12185_),
    .Y(_03753_));
 sky130_fd_sc_hd__o211a_1 _18919_ (.A1(_03222_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _18920_ (.A0(_03754_),
    .A1(net2445),
    .S(_03741_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _18921_ (.A(_03755_),
    .X(_00539_));
 sky130_fd_sc_hd__nand2_1 _18922_ (.A(_03752_),
    .B(_12198_),
    .Y(_03756_));
 sky130_fd_sc_hd__o211a_1 _18923_ (.A1(_03228_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__mux2_1 _18924_ (.A0(_03757_),
    .A1(net2607),
    .S(_03741_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _18925_ (.A(_03758_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _18926_ (.A(_03752_),
    .B(_12206_),
    .Y(_03759_));
 sky130_fd_sc_hd__o211a_1 _18927_ (.A1(_03232_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_1 _18928_ (.A0(_03760_),
    .A1(net2633),
    .S(_03741_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _18929_ (.A(_03761_),
    .X(_00541_));
 sky130_fd_sc_hd__nand2_1 _18930_ (.A(_03752_),
    .B(_12214_),
    .Y(_03762_));
 sky130_fd_sc_hd__o211a_1 _18931_ (.A1(_03236_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__mux2_1 _18932_ (.A0(_03763_),
    .A1(net2400),
    .S(_03741_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _18933_ (.A(_03764_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_1 _18934_ (.A(_03752_),
    .B(_12222_),
    .Y(_03765_));
 sky130_fd_sc_hd__o211a_1 _18935_ (.A1(_03240_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__mux2_1 _18936_ (.A0(_03766_),
    .A1(net2404),
    .S(_03741_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_1 _18937_ (.A(_03767_),
    .X(_00543_));
 sky130_fd_sc_hd__nand2_1 _18938_ (.A(_03752_),
    .B(_12230_),
    .Y(_03768_));
 sky130_fd_sc_hd__o211a_1 _18939_ (.A1(_03244_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_1 _18940_ (.A0(_03769_),
    .A1(net3307),
    .S(_03741_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _18941_ (.A(_03770_),
    .X(_00544_));
 sky130_fd_sc_hd__nand2_1 _18942_ (.A(_03752_),
    .B(_12238_),
    .Y(_03771_));
 sky130_fd_sc_hd__o211a_1 _18943_ (.A1(_03248_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__mux2_1 _18944_ (.A0(_03772_),
    .A1(net3515),
    .S(_03741_),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_1 _18945_ (.A(_03773_),
    .X(_00545_));
 sky130_fd_sc_hd__nand2_1 _18946_ (.A(_03752_),
    .B(_12246_),
    .Y(_03774_));
 sky130_fd_sc_hd__o211a_1 _18947_ (.A1(_03252_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__mux2_1 _18948_ (.A0(_03775_),
    .A1(net2533),
    .S(_03741_),
    .X(_03776_));
 sky130_fd_sc_hd__clkbuf_1 _18949_ (.A(_03776_),
    .X(_00546_));
 sky130_fd_sc_hd__o211a_1 _18950_ (.A1(_03256_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03753_),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_8 _18951_ (.A(_03740_),
    .X(_03778_));
 sky130_fd_sc_hd__mux2_1 _18952_ (.A0(_03777_),
    .A1(net3225),
    .S(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__clkbuf_1 _18953_ (.A(_03779_),
    .X(_00547_));
 sky130_fd_sc_hd__o211a_1 _18954_ (.A1(_03261_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03756_),
    .X(_03780_));
 sky130_fd_sc_hd__mux2_1 _18955_ (.A0(_03780_),
    .A1(net3420),
    .S(_03778_),
    .X(_03781_));
 sky130_fd_sc_hd__clkbuf_1 _18956_ (.A(_03781_),
    .X(_00548_));
 sky130_fd_sc_hd__o211a_1 _18957_ (.A1(_03264_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03759_),
    .X(_03782_));
 sky130_fd_sc_hd__mux2_1 _18958_ (.A0(_03782_),
    .A1(net2546),
    .S(_03778_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_1 _18959_ (.A(_03783_),
    .X(_00549_));
 sky130_fd_sc_hd__o211a_1 _18960_ (.A1(_03267_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03762_),
    .X(_03784_));
 sky130_fd_sc_hd__mux2_1 _18961_ (.A0(_03784_),
    .A1(net2448),
    .S(_03778_),
    .X(_03785_));
 sky130_fd_sc_hd__clkbuf_1 _18962_ (.A(_03785_),
    .X(_00550_));
 sky130_fd_sc_hd__o211a_1 _18963_ (.A1(_03270_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03765_),
    .X(_03786_));
 sky130_fd_sc_hd__mux2_1 _18964_ (.A0(_03786_),
    .A1(net3156),
    .S(_03778_),
    .X(_03787_));
 sky130_fd_sc_hd__clkbuf_1 _18965_ (.A(_03787_),
    .X(_00551_));
 sky130_fd_sc_hd__o211a_1 _18966_ (.A1(_03273_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03768_),
    .X(_03788_));
 sky130_fd_sc_hd__mux2_1 _18967_ (.A0(_03788_),
    .A1(net2416),
    .S(_03778_),
    .X(_03789_));
 sky130_fd_sc_hd__clkbuf_1 _18968_ (.A(_03789_),
    .X(_00552_));
 sky130_fd_sc_hd__o211a_1 _18969_ (.A1(_03276_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03771_),
    .X(_03790_));
 sky130_fd_sc_hd__mux2_1 _18970_ (.A0(_03790_),
    .A1(net2460),
    .S(_03778_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_1 _18971_ (.A(_03791_),
    .X(_00553_));
 sky130_fd_sc_hd__o211a_1 _18972_ (.A1(_03279_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03774_),
    .X(_03792_));
 sky130_fd_sc_hd__mux2_1 _18973_ (.A0(_03792_),
    .A1(net3135),
    .S(_03778_),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_1 _18974_ (.A(_03793_),
    .X(_00554_));
 sky130_fd_sc_hd__buf_4 _18975_ (.A(_03702_),
    .X(_03794_));
 sky130_fd_sc_hd__o211a_1 _18976_ (.A1(_12170_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03753_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _18977_ (.A0(_03795_),
    .A1(net3379),
    .S(_03778_),
    .X(_03796_));
 sky130_fd_sc_hd__clkbuf_1 _18978_ (.A(_03796_),
    .X(_00555_));
 sky130_fd_sc_hd__o211a_1 _18979_ (.A1(_12195_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03756_),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_1 _18980_ (.A0(_03797_),
    .A1(net2628),
    .S(_03778_),
    .X(_03798_));
 sky130_fd_sc_hd__clkbuf_1 _18981_ (.A(_03798_),
    .X(_00556_));
 sky130_fd_sc_hd__o211a_1 _18982_ (.A1(_12203_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03759_),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_1 _18983_ (.A0(_03799_),
    .A1(net3519),
    .S(_03778_),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_1 _18984_ (.A(_03800_),
    .X(_00557_));
 sky130_fd_sc_hd__o211a_1 _18985_ (.A1(_12211_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03762_),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _18986_ (.A0(_03801_),
    .A1(net3437),
    .S(_03778_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _18987_ (.A(_03802_),
    .X(_00558_));
 sky130_fd_sc_hd__o211a_1 _18988_ (.A1(_12219_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03765_),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_1 _18989_ (.A0(_03803_),
    .A1(net3689),
    .S(_03778_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_1 _18990_ (.A(_03804_),
    .X(_00559_));
 sky130_fd_sc_hd__o211a_1 _18991_ (.A1(_12227_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03768_),
    .X(_03805_));
 sky130_fd_sc_hd__mux2_1 _18992_ (.A0(_03805_),
    .A1(net3411),
    .S(_03778_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_1 _18993_ (.A(_03806_),
    .X(_00560_));
 sky130_fd_sc_hd__o211a_1 _18994_ (.A1(_12235_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03771_),
    .X(_03807_));
 sky130_fd_sc_hd__mux2_1 _18995_ (.A0(_03807_),
    .A1(net2461),
    .S(_03778_),
    .X(_03808_));
 sky130_fd_sc_hd__clkbuf_1 _18996_ (.A(_03808_),
    .X(_00561_));
 sky130_fd_sc_hd__o211a_1 _18997_ (.A1(_12243_),
    .A2(_03752_),
    .B1(_03794_),
    .C1(_03774_),
    .X(_03809_));
 sky130_fd_sc_hd__mux2_1 _18998_ (.A0(_03809_),
    .A1(net3679),
    .S(_03778_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _18999_ (.A(_03810_),
    .X(_00562_));
 sky130_fd_sc_hd__nor2_1 _19000_ (.A(_02812_),
    .B(_12175_),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2_2 _19001_ (.A(_03811_),
    .B(_12313_),
    .Y(_03812_));
 sky130_fd_sc_hd__buf_12 _19002_ (.A(_09109_),
    .X(_03813_));
 sky130_fd_sc_hd__a21bo_1 _19003_ (.A1(_03812_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_8 _19004_ (.A(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__mux2_1 _19005_ (.A0(_02810_),
    .A1(net2152),
    .S(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _19006_ (.A(_03816_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _19007_ (.A0(_02823_),
    .A1(net2198),
    .S(_03815_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_1 _19008_ (.A(_03817_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _19009_ (.A0(_02827_),
    .A1(net2189),
    .S(_03815_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _19010_ (.A(_03818_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _19011_ (.A0(_02831_),
    .A1(net3099),
    .S(_03815_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _19012_ (.A(_03819_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _19013_ (.A0(_02835_),
    .A1(net3231),
    .S(_03815_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _19014_ (.A(_03820_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _19015_ (.A0(_02839_),
    .A1(net2982),
    .S(_03815_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_1 _19016_ (.A(_03821_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _19017_ (.A0(_02843_),
    .A1(net2262),
    .S(_03815_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _19018_ (.A(_03822_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _19019_ (.A0(_02847_),
    .A1(net3604),
    .S(_03815_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _19020_ (.A(_03823_),
    .X(_00570_));
 sky130_fd_sc_hd__buf_4 _19021_ (.A(_03812_),
    .X(_03824_));
 sky130_fd_sc_hd__buf_4 _19022_ (.A(_03812_),
    .X(_03825_));
 sky130_fd_sc_hd__nand2_1 _19023_ (.A(_03825_),
    .B(_12185_),
    .Y(_03826_));
 sky130_fd_sc_hd__o211a_1 _19024_ (.A1(_03222_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__mux2_1 _19025_ (.A0(_03827_),
    .A1(net2388),
    .S(_03815_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_1 _19026_ (.A(_03828_),
    .X(_00571_));
 sky130_fd_sc_hd__nand2_1 _19027_ (.A(_03825_),
    .B(_12198_),
    .Y(_03829_));
 sky130_fd_sc_hd__o211a_1 _19028_ (.A1(_03228_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _19029_ (.A0(_03830_),
    .A1(net3086),
    .S(_03815_),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _19030_ (.A(_03831_),
    .X(_00572_));
 sky130_fd_sc_hd__nand2_1 _19031_ (.A(_03825_),
    .B(_12206_),
    .Y(_03832_));
 sky130_fd_sc_hd__o211a_1 _19032_ (.A1(_03232_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__mux2_1 _19033_ (.A0(_03833_),
    .A1(net2383),
    .S(_03815_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _19034_ (.A(_03834_),
    .X(_00573_));
 sky130_fd_sc_hd__nand2_1 _19035_ (.A(_03825_),
    .B(_12214_),
    .Y(_03835_));
 sky130_fd_sc_hd__o211a_1 _19036_ (.A1(_03236_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_1 _19037_ (.A0(_03836_),
    .A1(net2843),
    .S(_03815_),
    .X(_03837_));
 sky130_fd_sc_hd__clkbuf_1 _19038_ (.A(_03837_),
    .X(_00574_));
 sky130_fd_sc_hd__nand2_1 _19039_ (.A(_03825_),
    .B(_12222_),
    .Y(_03838_));
 sky130_fd_sc_hd__o211a_1 _19040_ (.A1(_03240_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _19041_ (.A0(_03839_),
    .A1(net2946),
    .S(_03815_),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_1 _19042_ (.A(_03840_),
    .X(_00575_));
 sky130_fd_sc_hd__nand2_1 _19043_ (.A(_03825_),
    .B(_12230_),
    .Y(_03841_));
 sky130_fd_sc_hd__o211a_1 _19044_ (.A1(_03244_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__mux2_1 _19045_ (.A0(_03842_),
    .A1(net2783),
    .S(_03815_),
    .X(_03843_));
 sky130_fd_sc_hd__clkbuf_1 _19046_ (.A(_03843_),
    .X(_00576_));
 sky130_fd_sc_hd__nand2_1 _19047_ (.A(_03825_),
    .B(_12238_),
    .Y(_03844_));
 sky130_fd_sc_hd__o211a_1 _19048_ (.A1(_03248_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__mux2_1 _19049_ (.A0(_03845_),
    .A1(net2303),
    .S(_03815_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _19050_ (.A(_03846_),
    .X(_00577_));
 sky130_fd_sc_hd__nand2_1 _19051_ (.A(_03825_),
    .B(_12246_),
    .Y(_03847_));
 sky130_fd_sc_hd__o211a_1 _19052_ (.A1(_03252_),
    .A2(_03824_),
    .B1(_03794_),
    .C1(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__mux2_1 _19053_ (.A0(_03848_),
    .A1(net3100),
    .S(_03815_),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_1 _19054_ (.A(_03849_),
    .X(_00578_));
 sky130_fd_sc_hd__buf_4 _19055_ (.A(_03702_),
    .X(_03850_));
 sky130_fd_sc_hd__o211a_1 _19056_ (.A1(_03256_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03826_),
    .X(_03851_));
 sky130_fd_sc_hd__clkbuf_8 _19057_ (.A(_03814_),
    .X(_03852_));
 sky130_fd_sc_hd__mux2_1 _19058_ (.A0(_03851_),
    .A1(net3051),
    .S(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_1 _19059_ (.A(_03853_),
    .X(_00579_));
 sky130_fd_sc_hd__o211a_1 _19060_ (.A1(_03261_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03829_),
    .X(_03854_));
 sky130_fd_sc_hd__mux2_1 _19061_ (.A0(_03854_),
    .A1(net2473),
    .S(_03852_),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_1 _19062_ (.A(_03855_),
    .X(_00580_));
 sky130_fd_sc_hd__o211a_1 _19063_ (.A1(_03264_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03832_),
    .X(_03856_));
 sky130_fd_sc_hd__mux2_1 _19064_ (.A0(_03856_),
    .A1(net2406),
    .S(_03852_),
    .X(_03857_));
 sky130_fd_sc_hd__clkbuf_1 _19065_ (.A(_03857_),
    .X(_00581_));
 sky130_fd_sc_hd__o211a_1 _19066_ (.A1(_03267_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03835_),
    .X(_03858_));
 sky130_fd_sc_hd__mux2_1 _19067_ (.A0(_03858_),
    .A1(net3525),
    .S(_03852_),
    .X(_03859_));
 sky130_fd_sc_hd__clkbuf_1 _19068_ (.A(_03859_),
    .X(_00582_));
 sky130_fd_sc_hd__o211a_1 _19069_ (.A1(_03270_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03838_),
    .X(_03860_));
 sky130_fd_sc_hd__mux2_1 _19070_ (.A0(_03860_),
    .A1(net2816),
    .S(_03852_),
    .X(_03861_));
 sky130_fd_sc_hd__clkbuf_1 _19071_ (.A(_03861_),
    .X(_00583_));
 sky130_fd_sc_hd__o211a_1 _19072_ (.A1(_03273_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03841_),
    .X(_03862_));
 sky130_fd_sc_hd__mux2_1 _19073_ (.A0(_03862_),
    .A1(net2456),
    .S(_03852_),
    .X(_03863_));
 sky130_fd_sc_hd__clkbuf_1 _19074_ (.A(_03863_),
    .X(_00584_));
 sky130_fd_sc_hd__o211a_1 _19075_ (.A1(_03276_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03844_),
    .X(_03864_));
 sky130_fd_sc_hd__mux2_1 _19076_ (.A0(_03864_),
    .A1(net2662),
    .S(_03852_),
    .X(_03865_));
 sky130_fd_sc_hd__clkbuf_1 _19077_ (.A(_03865_),
    .X(_00585_));
 sky130_fd_sc_hd__o211a_1 _19078_ (.A1(_03279_),
    .A2(_03824_),
    .B1(_03850_),
    .C1(_03847_),
    .X(_03866_));
 sky130_fd_sc_hd__mux2_1 _19079_ (.A0(_03866_),
    .A1(net2720),
    .S(_03852_),
    .X(_03867_));
 sky130_fd_sc_hd__clkbuf_1 _19080_ (.A(_03867_),
    .X(_00586_));
 sky130_fd_sc_hd__o211a_1 _19081_ (.A1(_12170_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03826_),
    .X(_03868_));
 sky130_fd_sc_hd__mux2_1 _19082_ (.A0(_03868_),
    .A1(net3141),
    .S(_03852_),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_1 _19083_ (.A(_03869_),
    .X(_00587_));
 sky130_fd_sc_hd__o211a_1 _19084_ (.A1(_12195_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03829_),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _19085_ (.A0(_03870_),
    .A1(net2171),
    .S(_03852_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _19086_ (.A(_03871_),
    .X(_00588_));
 sky130_fd_sc_hd__o211a_1 _19087_ (.A1(_12203_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03832_),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _19088_ (.A0(_03872_),
    .A1(net2246),
    .S(_03852_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _19089_ (.A(_03873_),
    .X(_00589_));
 sky130_fd_sc_hd__o211a_1 _19090_ (.A1(_12211_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03835_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _19091_ (.A0(_03874_),
    .A1(net2538),
    .S(_03852_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_1 _19092_ (.A(_03875_),
    .X(_00590_));
 sky130_fd_sc_hd__o211a_1 _19093_ (.A1(_12219_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03838_),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _19094_ (.A0(_03876_),
    .A1(net2700),
    .S(_03852_),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_1 _19095_ (.A(_03877_),
    .X(_00591_));
 sky130_fd_sc_hd__o211a_1 _19096_ (.A1(_12227_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03841_),
    .X(_03878_));
 sky130_fd_sc_hd__mux2_1 _19097_ (.A0(_03878_),
    .A1(net2414),
    .S(_03852_),
    .X(_03879_));
 sky130_fd_sc_hd__clkbuf_1 _19098_ (.A(_03879_),
    .X(_00592_));
 sky130_fd_sc_hd__o211a_1 _19099_ (.A1(_12235_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03844_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_1 _19100_ (.A0(_03880_),
    .A1(net2651),
    .S(_03852_),
    .X(_03881_));
 sky130_fd_sc_hd__clkbuf_1 _19101_ (.A(_03881_),
    .X(_00593_));
 sky130_fd_sc_hd__o211a_1 _19102_ (.A1(_12243_),
    .A2(_03825_),
    .B1(_03850_),
    .C1(_03847_),
    .X(_03882_));
 sky130_fd_sc_hd__mux2_1 _19103_ (.A0(_03882_),
    .A1(net3253),
    .S(_03852_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_1 _19104_ (.A(_03883_),
    .X(_00594_));
 sky130_fd_sc_hd__nor2_1 _19105_ (.A(_12293_),
    .B(_12175_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_2 _19106_ (.A(_03884_),
    .B(_12313_),
    .Y(_03885_));
 sky130_fd_sc_hd__a21bo_1 _19107_ (.A1(_03885_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_03886_));
 sky130_fd_sc_hd__clkbuf_8 _19108_ (.A(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__mux2_1 _19109_ (.A0(_02810_),
    .A1(net3128),
    .S(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__clkbuf_1 _19110_ (.A(_03888_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _19111_ (.A0(_02823_),
    .A1(net3351),
    .S(_03887_),
    .X(_03889_));
 sky130_fd_sc_hd__clkbuf_1 _19112_ (.A(_03889_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _19113_ (.A0(_02827_),
    .A1(net3283),
    .S(_03887_),
    .X(_03890_));
 sky130_fd_sc_hd__clkbuf_1 _19114_ (.A(_03890_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _19115_ (.A0(_02831_),
    .A1(net3334),
    .S(_03887_),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_1 _19116_ (.A(_03891_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _19117_ (.A0(_02835_),
    .A1(net2966),
    .S(_03887_),
    .X(_03892_));
 sky130_fd_sc_hd__clkbuf_1 _19118_ (.A(_03892_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _19119_ (.A0(_02839_),
    .A1(net3230),
    .S(_03887_),
    .X(_03893_));
 sky130_fd_sc_hd__clkbuf_1 _19120_ (.A(_03893_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _19121_ (.A0(_02843_),
    .A1(net2492),
    .S(_03887_),
    .X(_03894_));
 sky130_fd_sc_hd__clkbuf_1 _19122_ (.A(_03894_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _19123_ (.A0(_02847_),
    .A1(net2858),
    .S(_03887_),
    .X(_03895_));
 sky130_fd_sc_hd__clkbuf_1 _19124_ (.A(_03895_),
    .X(_00602_));
 sky130_fd_sc_hd__buf_4 _19125_ (.A(_03885_),
    .X(_03896_));
 sky130_fd_sc_hd__buf_4 _19126_ (.A(_03702_),
    .X(_03897_));
 sky130_fd_sc_hd__buf_4 _19127_ (.A(_03885_),
    .X(_03898_));
 sky130_fd_sc_hd__nand2_1 _19128_ (.A(_03898_),
    .B(_12185_),
    .Y(_03899_));
 sky130_fd_sc_hd__o211a_1 _19129_ (.A1(_03222_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_1 _19130_ (.A0(_03900_),
    .A1(net2707),
    .S(_03887_),
    .X(_03901_));
 sky130_fd_sc_hd__clkbuf_1 _19131_ (.A(_03901_),
    .X(_00603_));
 sky130_fd_sc_hd__nand2_1 _19132_ (.A(_03898_),
    .B(_12198_),
    .Y(_03902_));
 sky130_fd_sc_hd__o211a_1 _19133_ (.A1(_03228_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__mux2_1 _19134_ (.A0(_03903_),
    .A1(net2300),
    .S(_03887_),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_1 _19135_ (.A(_03904_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _19136_ (.A(_03898_),
    .B(_12206_),
    .Y(_03905_));
 sky130_fd_sc_hd__o211a_1 _19137_ (.A1(_03232_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__mux2_1 _19138_ (.A0(_03906_),
    .A1(net3298),
    .S(_03887_),
    .X(_03907_));
 sky130_fd_sc_hd__clkbuf_1 _19139_ (.A(_03907_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _19140_ (.A(_03898_),
    .B(_12214_),
    .Y(_03908_));
 sky130_fd_sc_hd__o211a_1 _19141_ (.A1(_03236_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _19142_ (.A0(_03909_),
    .A1(net3214),
    .S(_03887_),
    .X(_03910_));
 sky130_fd_sc_hd__clkbuf_1 _19143_ (.A(_03910_),
    .X(_00606_));
 sky130_fd_sc_hd__nand2_1 _19144_ (.A(_03898_),
    .B(_12222_),
    .Y(_03911_));
 sky130_fd_sc_hd__o211a_1 _19145_ (.A1(_03240_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__mux2_1 _19146_ (.A0(_03912_),
    .A1(net2894),
    .S(_03887_),
    .X(_03913_));
 sky130_fd_sc_hd__clkbuf_1 _19147_ (.A(_03913_),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _19148_ (.A(_03898_),
    .B(_12230_),
    .Y(_03914_));
 sky130_fd_sc_hd__o211a_1 _19149_ (.A1(_03244_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_1 _19150_ (.A0(_03915_),
    .A1(net3258),
    .S(_03887_),
    .X(_03916_));
 sky130_fd_sc_hd__clkbuf_1 _19151_ (.A(_03916_),
    .X(_00608_));
 sky130_fd_sc_hd__nand2_1 _19152_ (.A(_03898_),
    .B(_12238_),
    .Y(_03917_));
 sky130_fd_sc_hd__o211a_1 _19153_ (.A1(_03248_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_1 _19154_ (.A0(_03918_),
    .A1(net3180),
    .S(_03887_),
    .X(_03919_));
 sky130_fd_sc_hd__clkbuf_1 _19155_ (.A(_03919_),
    .X(_00609_));
 sky130_fd_sc_hd__nand2_1 _19156_ (.A(_03898_),
    .B(_12246_),
    .Y(_03920_));
 sky130_fd_sc_hd__o211a_1 _19157_ (.A1(_03252_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_1 _19158_ (.A0(_03921_),
    .A1(net2398),
    .S(_03887_),
    .X(_03922_));
 sky130_fd_sc_hd__clkbuf_1 _19159_ (.A(_03922_),
    .X(_00610_));
 sky130_fd_sc_hd__o211a_1 _19160_ (.A1(_03256_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03899_),
    .X(_03923_));
 sky130_fd_sc_hd__clkbuf_8 _19161_ (.A(_03886_),
    .X(_03924_));
 sky130_fd_sc_hd__mux2_1 _19162_ (.A0(_03923_),
    .A1(net2376),
    .S(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__clkbuf_1 _19163_ (.A(_03925_),
    .X(_00611_));
 sky130_fd_sc_hd__o211a_1 _19164_ (.A1(_03261_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03902_),
    .X(_03926_));
 sky130_fd_sc_hd__mux2_1 _19165_ (.A0(_03926_),
    .A1(net2933),
    .S(_03924_),
    .X(_03927_));
 sky130_fd_sc_hd__clkbuf_1 _19166_ (.A(_03927_),
    .X(_00612_));
 sky130_fd_sc_hd__o211a_1 _19167_ (.A1(_03264_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03905_),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_1 _19168_ (.A0(_03928_),
    .A1(net3200),
    .S(_03924_),
    .X(_03929_));
 sky130_fd_sc_hd__clkbuf_1 _19169_ (.A(_03929_),
    .X(_00613_));
 sky130_fd_sc_hd__o211a_1 _19170_ (.A1(_03267_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03908_),
    .X(_03930_));
 sky130_fd_sc_hd__mux2_1 _19171_ (.A0(_03930_),
    .A1(net3157),
    .S(_03924_),
    .X(_03931_));
 sky130_fd_sc_hd__clkbuf_1 _19172_ (.A(_03931_),
    .X(_00614_));
 sky130_fd_sc_hd__o211a_1 _19173_ (.A1(_03270_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03911_),
    .X(_03932_));
 sky130_fd_sc_hd__mux2_1 _19174_ (.A0(_03932_),
    .A1(net3339),
    .S(_03924_),
    .X(_03933_));
 sky130_fd_sc_hd__clkbuf_1 _19175_ (.A(_03933_),
    .X(_00615_));
 sky130_fd_sc_hd__o211a_1 _19176_ (.A1(_03273_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03914_),
    .X(_03934_));
 sky130_fd_sc_hd__mux2_1 _19177_ (.A0(_03934_),
    .A1(net3149),
    .S(_03924_),
    .X(_03935_));
 sky130_fd_sc_hd__clkbuf_1 _19178_ (.A(_03935_),
    .X(_00616_));
 sky130_fd_sc_hd__o211a_1 _19179_ (.A1(_03276_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03917_),
    .X(_03936_));
 sky130_fd_sc_hd__mux2_1 _19180_ (.A0(_03936_),
    .A1(net2953),
    .S(_03924_),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_1 _19181_ (.A(_03937_),
    .X(_00617_));
 sky130_fd_sc_hd__o211a_1 _19182_ (.A1(_03279_),
    .A2(_03896_),
    .B1(_03897_),
    .C1(_03920_),
    .X(_03938_));
 sky130_fd_sc_hd__mux2_1 _19183_ (.A0(_03938_),
    .A1(net2496),
    .S(_03924_),
    .X(_03939_));
 sky130_fd_sc_hd__clkbuf_1 _19184_ (.A(_03939_),
    .X(_00618_));
 sky130_fd_sc_hd__buf_4 _19185_ (.A(_03702_),
    .X(_03940_));
 sky130_fd_sc_hd__o211a_1 _19186_ (.A1(_12170_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03899_),
    .X(_03941_));
 sky130_fd_sc_hd__mux2_1 _19187_ (.A0(_03941_),
    .A1(net2588),
    .S(_03924_),
    .X(_03942_));
 sky130_fd_sc_hd__clkbuf_1 _19188_ (.A(_03942_),
    .X(_00619_));
 sky130_fd_sc_hd__o211a_1 _19189_ (.A1(_12195_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03902_),
    .X(_03943_));
 sky130_fd_sc_hd__mux2_1 _19190_ (.A0(_03943_),
    .A1(net3505),
    .S(_03924_),
    .X(_03944_));
 sky130_fd_sc_hd__clkbuf_1 _19191_ (.A(_03944_),
    .X(_00620_));
 sky130_fd_sc_hd__o211a_1 _19192_ (.A1(_12203_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03905_),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_1 _19193_ (.A0(_03945_),
    .A1(net3039),
    .S(_03924_),
    .X(_03946_));
 sky130_fd_sc_hd__clkbuf_1 _19194_ (.A(_03946_),
    .X(_00621_));
 sky130_fd_sc_hd__o211a_1 _19195_ (.A1(_12211_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03908_),
    .X(_03947_));
 sky130_fd_sc_hd__mux2_1 _19196_ (.A0(_03947_),
    .A1(net2614),
    .S(_03924_),
    .X(_03948_));
 sky130_fd_sc_hd__clkbuf_1 _19197_ (.A(_03948_),
    .X(_00622_));
 sky130_fd_sc_hd__o211a_1 _19198_ (.A1(_12219_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03911_),
    .X(_03949_));
 sky130_fd_sc_hd__mux2_1 _19199_ (.A0(_03949_),
    .A1(net3207),
    .S(_03924_),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_1 _19200_ (.A(_03950_),
    .X(_00623_));
 sky130_fd_sc_hd__o211a_1 _19201_ (.A1(_12227_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03914_),
    .X(_03951_));
 sky130_fd_sc_hd__mux2_1 _19202_ (.A0(_03951_),
    .A1(net3001),
    .S(_03924_),
    .X(_03952_));
 sky130_fd_sc_hd__clkbuf_1 _19203_ (.A(_03952_),
    .X(_00624_));
 sky130_fd_sc_hd__o211a_1 _19204_ (.A1(_12235_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03917_),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_1 _19205_ (.A0(_03953_),
    .A1(net2897),
    .S(_03924_),
    .X(_03954_));
 sky130_fd_sc_hd__clkbuf_1 _19206_ (.A(_03954_),
    .X(_00625_));
 sky130_fd_sc_hd__o211a_1 _19207_ (.A1(_12243_),
    .A2(_03898_),
    .B1(_03940_),
    .C1(_03920_),
    .X(_03955_));
 sky130_fd_sc_hd__mux2_1 _19208_ (.A0(_03955_),
    .A1(net3355),
    .S(_03924_),
    .X(_03956_));
 sky130_fd_sc_hd__clkbuf_1 _19209_ (.A(_03956_),
    .X(_00626_));
 sky130_fd_sc_hd__nor2_1 _19210_ (.A(_12292_),
    .B(_12175_),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2_2 _19211_ (.A(_03957_),
    .B(_12313_),
    .Y(_03958_));
 sky130_fd_sc_hd__a21bo_1 _19212_ (.A1(_03958_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_03959_));
 sky130_fd_sc_hd__clkbuf_8 _19213_ (.A(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__mux2_1 _19214_ (.A0(_02810_),
    .A1(net2873),
    .S(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__clkbuf_1 _19215_ (.A(_03961_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _19216_ (.A0(_02823_),
    .A1(net2255),
    .S(_03960_),
    .X(_03962_));
 sky130_fd_sc_hd__clkbuf_1 _19217_ (.A(_03962_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _19218_ (.A0(_02827_),
    .A1(net2744),
    .S(_03960_),
    .X(_03963_));
 sky130_fd_sc_hd__clkbuf_1 _19219_ (.A(_03963_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _19220_ (.A0(_02831_),
    .A1(net2326),
    .S(_03960_),
    .X(_03964_));
 sky130_fd_sc_hd__clkbuf_1 _19221_ (.A(_03964_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _19222_ (.A0(_02835_),
    .A1(net2267),
    .S(_03960_),
    .X(_03965_));
 sky130_fd_sc_hd__clkbuf_1 _19223_ (.A(_03965_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _19224_ (.A0(_02839_),
    .A1(net2494),
    .S(_03960_),
    .X(_03966_));
 sky130_fd_sc_hd__clkbuf_1 _19225_ (.A(_03966_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _19226_ (.A0(_02843_),
    .A1(net2769),
    .S(_03960_),
    .X(_03967_));
 sky130_fd_sc_hd__clkbuf_1 _19227_ (.A(_03967_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _19228_ (.A0(_02847_),
    .A1(net2149),
    .S(_03960_),
    .X(_03968_));
 sky130_fd_sc_hd__clkbuf_1 _19229_ (.A(_03968_),
    .X(_00634_));
 sky130_fd_sc_hd__buf_4 _19230_ (.A(_03958_),
    .X(_03969_));
 sky130_fd_sc_hd__buf_4 _19231_ (.A(_03958_),
    .X(_03970_));
 sky130_fd_sc_hd__nand2_1 _19232_ (.A(_03970_),
    .B(_12185_),
    .Y(_03971_));
 sky130_fd_sc_hd__o211a_1 _19233_ (.A1(_03222_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__mux2_1 _19234_ (.A0(_03972_),
    .A1(net3343),
    .S(_03960_),
    .X(_03973_));
 sky130_fd_sc_hd__clkbuf_1 _19235_ (.A(_03973_),
    .X(_00635_));
 sky130_fd_sc_hd__nand2_1 _19236_ (.A(_03970_),
    .B(_12198_),
    .Y(_03974_));
 sky130_fd_sc_hd__o211a_1 _19237_ (.A1(_03228_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _19238_ (.A0(_03975_),
    .A1(net3588),
    .S(_03960_),
    .X(_03976_));
 sky130_fd_sc_hd__clkbuf_1 _19239_ (.A(_03976_),
    .X(_00636_));
 sky130_fd_sc_hd__nand2_1 _19240_ (.A(_03970_),
    .B(_12206_),
    .Y(_03977_));
 sky130_fd_sc_hd__o211a_1 _19241_ (.A1(_03232_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__mux2_1 _19242_ (.A0(_03978_),
    .A1(net3480),
    .S(_03960_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_1 _19243_ (.A(_03979_),
    .X(_00637_));
 sky130_fd_sc_hd__nand2_1 _19244_ (.A(_03970_),
    .B(_12214_),
    .Y(_03980_));
 sky130_fd_sc_hd__o211a_1 _19245_ (.A1(_03236_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__mux2_1 _19246_ (.A0(_03981_),
    .A1(net3144),
    .S(_03960_),
    .X(_03982_));
 sky130_fd_sc_hd__clkbuf_1 _19247_ (.A(_03982_),
    .X(_00638_));
 sky130_fd_sc_hd__nand2_1 _19248_ (.A(_03970_),
    .B(_12222_),
    .Y(_03983_));
 sky130_fd_sc_hd__o211a_1 _19249_ (.A1(_03240_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__mux2_1 _19250_ (.A0(_03984_),
    .A1(net3315),
    .S(_03960_),
    .X(_03985_));
 sky130_fd_sc_hd__clkbuf_1 _19251_ (.A(_03985_),
    .X(_00639_));
 sky130_fd_sc_hd__nand2_1 _19252_ (.A(_03970_),
    .B(_12230_),
    .Y(_03986_));
 sky130_fd_sc_hd__o211a_1 _19253_ (.A1(_03244_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_1 _19254_ (.A0(_03987_),
    .A1(net3020),
    .S(_03960_),
    .X(_03988_));
 sky130_fd_sc_hd__clkbuf_1 _19255_ (.A(_03988_),
    .X(_00640_));
 sky130_fd_sc_hd__nand2_1 _19256_ (.A(_03970_),
    .B(_12238_),
    .Y(_03989_));
 sky130_fd_sc_hd__o211a_1 _19257_ (.A1(_03248_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__mux2_1 _19258_ (.A0(_03990_),
    .A1(net3582),
    .S(_03960_),
    .X(_03991_));
 sky130_fd_sc_hd__clkbuf_1 _19259_ (.A(_03991_),
    .X(_00641_));
 sky130_fd_sc_hd__nand2_1 _19260_ (.A(_03970_),
    .B(_12246_),
    .Y(_03992_));
 sky130_fd_sc_hd__o211a_1 _19261_ (.A1(_03252_),
    .A2(_03969_),
    .B1(_03940_),
    .C1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _19262_ (.A0(_03993_),
    .A1(net3360),
    .S(_03960_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_1 _19263_ (.A(_03994_),
    .X(_00642_));
 sky130_fd_sc_hd__buf_4 _19264_ (.A(_03702_),
    .X(_03995_));
 sky130_fd_sc_hd__o211a_1 _19265_ (.A1(_03256_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03971_),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_8 _19266_ (.A(_03959_),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_1 _19267_ (.A0(_03996_),
    .A1(net3204),
    .S(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__clkbuf_1 _19268_ (.A(_03998_),
    .X(_00643_));
 sky130_fd_sc_hd__o211a_1 _19269_ (.A1(_03261_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03974_),
    .X(_03999_));
 sky130_fd_sc_hd__mux2_1 _19270_ (.A0(_03999_),
    .A1(net3371),
    .S(_03997_),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_1 _19271_ (.A(_04000_),
    .X(_00644_));
 sky130_fd_sc_hd__o211a_1 _19272_ (.A1(_03264_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03977_),
    .X(_04001_));
 sky130_fd_sc_hd__mux2_1 _19273_ (.A0(_04001_),
    .A1(net3537),
    .S(_03997_),
    .X(_04002_));
 sky130_fd_sc_hd__clkbuf_1 _19274_ (.A(_04002_),
    .X(_00645_));
 sky130_fd_sc_hd__o211a_1 _19275_ (.A1(_03267_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03980_),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_1 _19276_ (.A0(_04003_),
    .A1(net3650),
    .S(_03997_),
    .X(_04004_));
 sky130_fd_sc_hd__clkbuf_1 _19277_ (.A(_04004_),
    .X(_00646_));
 sky130_fd_sc_hd__o211a_1 _19278_ (.A1(_03270_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03983_),
    .X(_04005_));
 sky130_fd_sc_hd__mux2_1 _19279_ (.A0(_04005_),
    .A1(net2215),
    .S(_03997_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_1 _19280_ (.A(_04006_),
    .X(_00647_));
 sky130_fd_sc_hd__o211a_1 _19281_ (.A1(_03273_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03986_),
    .X(_04007_));
 sky130_fd_sc_hd__mux2_1 _19282_ (.A0(_04007_),
    .A1(net2755),
    .S(_03997_),
    .X(_04008_));
 sky130_fd_sc_hd__clkbuf_1 _19283_ (.A(_04008_),
    .X(_00648_));
 sky130_fd_sc_hd__o211a_1 _19284_ (.A1(_03276_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03989_),
    .X(_04009_));
 sky130_fd_sc_hd__mux2_1 _19285_ (.A0(_04009_),
    .A1(net3304),
    .S(_03997_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_1 _19286_ (.A(_04010_),
    .X(_00649_));
 sky130_fd_sc_hd__o211a_1 _19287_ (.A1(_03279_),
    .A2(_03969_),
    .B1(_03995_),
    .C1(_03992_),
    .X(_04011_));
 sky130_fd_sc_hd__mux2_1 _19288_ (.A0(_04011_),
    .A1(net3038),
    .S(_03997_),
    .X(_04012_));
 sky130_fd_sc_hd__clkbuf_1 _19289_ (.A(_04012_),
    .X(_00650_));
 sky130_fd_sc_hd__o211a_1 _19290_ (.A1(_12170_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03971_),
    .X(_04013_));
 sky130_fd_sc_hd__mux2_1 _19291_ (.A0(_04013_),
    .A1(net2446),
    .S(_03997_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _19292_ (.A(_04014_),
    .X(_00651_));
 sky130_fd_sc_hd__o211a_1 _19293_ (.A1(_12195_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03974_),
    .X(_04015_));
 sky130_fd_sc_hd__mux2_1 _19294_ (.A0(_04015_),
    .A1(net3700),
    .S(_03997_),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_1 _19295_ (.A(_04016_),
    .X(_00652_));
 sky130_fd_sc_hd__o211a_1 _19296_ (.A1(_12203_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03977_),
    .X(_04017_));
 sky130_fd_sc_hd__mux2_1 _19297_ (.A0(_04017_),
    .A1(net3391),
    .S(_03997_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _19298_ (.A(_04018_),
    .X(_00653_));
 sky130_fd_sc_hd__o211a_1 _19299_ (.A1(_12211_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03980_),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _19300_ (.A0(_04019_),
    .A1(net2594),
    .S(_03997_),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_1 _19301_ (.A(_04020_),
    .X(_00654_));
 sky130_fd_sc_hd__o211a_1 _19302_ (.A1(_12219_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03983_),
    .X(_04021_));
 sky130_fd_sc_hd__mux2_1 _19303_ (.A0(_04021_),
    .A1(net2997),
    .S(_03997_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _19304_ (.A(_04022_),
    .X(_00655_));
 sky130_fd_sc_hd__o211a_1 _19305_ (.A1(_12227_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03986_),
    .X(_04023_));
 sky130_fd_sc_hd__mux2_1 _19306_ (.A0(_04023_),
    .A1(net2213),
    .S(_03997_),
    .X(_04024_));
 sky130_fd_sc_hd__clkbuf_1 _19307_ (.A(_04024_),
    .X(_00656_));
 sky130_fd_sc_hd__o211a_1 _19308_ (.A1(_12235_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03989_),
    .X(_04025_));
 sky130_fd_sc_hd__mux2_1 _19309_ (.A0(_04025_),
    .A1(net2314),
    .S(_03997_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_1 _19310_ (.A(_04026_),
    .X(_00657_));
 sky130_fd_sc_hd__o211a_1 _19311_ (.A1(_12243_),
    .A2(_03970_),
    .B1(_03995_),
    .C1(_03992_),
    .X(_04027_));
 sky130_fd_sc_hd__mux2_1 _19312_ (.A0(_04027_),
    .A1(net2931),
    .S(_03997_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _19313_ (.A(_04028_),
    .X(_00658_));
 sky130_fd_sc_hd__nand2_2 _19314_ (.A(_12176_),
    .B(_12313_),
    .Y(_04029_));
 sky130_fd_sc_hd__a21bo_1 _19315_ (.A1(_04029_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_04030_));
 sky130_fd_sc_hd__clkbuf_8 _19316_ (.A(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__mux2_1 _19317_ (.A0(_02810_),
    .A1(net2882),
    .S(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__clkbuf_1 _19318_ (.A(_04032_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _19319_ (.A0(_02823_),
    .A1(net2573),
    .S(_04031_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_1 _19320_ (.A(_04033_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _19321_ (.A0(_02827_),
    .A1(net2836),
    .S(_04031_),
    .X(_04034_));
 sky130_fd_sc_hd__clkbuf_1 _19322_ (.A(_04034_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _19323_ (.A0(_02831_),
    .A1(net2352),
    .S(_04031_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_1 _19324_ (.A(_04035_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _19325_ (.A0(_02835_),
    .A1(net3007),
    .S(_04031_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _19326_ (.A(_04036_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _19327_ (.A0(_02839_),
    .A1(net2577),
    .S(_04031_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _19328_ (.A(_04037_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _19329_ (.A0(_02843_),
    .A1(net3046),
    .S(_04031_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _19330_ (.A(_04038_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _19331_ (.A0(_02847_),
    .A1(net3003),
    .S(_04031_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_1 _19332_ (.A(_04039_),
    .X(_00666_));
 sky130_fd_sc_hd__buf_4 _19333_ (.A(_04029_),
    .X(_04040_));
 sky130_fd_sc_hd__buf_4 _19334_ (.A(_03702_),
    .X(_04041_));
 sky130_fd_sc_hd__buf_4 _19335_ (.A(_04029_),
    .X(_04042_));
 sky130_fd_sc_hd__nand2_1 _19336_ (.A(_04042_),
    .B(_12185_),
    .Y(_04043_));
 sky130_fd_sc_hd__o211a_1 _19337_ (.A1(_03222_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__mux2_1 _19338_ (.A0(_04044_),
    .A1(net3155),
    .S(_04031_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _19339_ (.A(_04045_),
    .X(_00667_));
 sky130_fd_sc_hd__nand2_1 _19340_ (.A(_04042_),
    .B(_12198_),
    .Y(_04046_));
 sky130_fd_sc_hd__o211a_1 _19341_ (.A1(_03228_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__mux2_1 _19342_ (.A0(_04047_),
    .A1(net2237),
    .S(_04031_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _19343_ (.A(_04048_),
    .X(_00668_));
 sky130_fd_sc_hd__nand2_1 _19344_ (.A(_04042_),
    .B(_12206_),
    .Y(_04049_));
 sky130_fd_sc_hd__o211a_1 _19345_ (.A1(_03232_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__mux2_1 _19346_ (.A0(_04050_),
    .A1(net2752),
    .S(_04031_),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_1 _19347_ (.A(_04051_),
    .X(_00669_));
 sky130_fd_sc_hd__nand2_1 _19348_ (.A(_04042_),
    .B(_12214_),
    .Y(_04052_));
 sky130_fd_sc_hd__o211a_1 _19349_ (.A1(_03236_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__mux2_1 _19350_ (.A0(_04053_),
    .A1(net2703),
    .S(_04031_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_1 _19351_ (.A(_04054_),
    .X(_00670_));
 sky130_fd_sc_hd__nand2_1 _19352_ (.A(_04042_),
    .B(_12222_),
    .Y(_04055_));
 sky130_fd_sc_hd__o211a_1 _19353_ (.A1(_03240_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__mux2_1 _19354_ (.A0(_04056_),
    .A1(net3446),
    .S(_04031_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _19355_ (.A(_04057_),
    .X(_00671_));
 sky130_fd_sc_hd__nand2_1 _19356_ (.A(_04042_),
    .B(_12230_),
    .Y(_04058_));
 sky130_fd_sc_hd__o211a_1 _19357_ (.A1(_03244_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__mux2_1 _19358_ (.A0(_04059_),
    .A1(net3601),
    .S(_04031_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _19359_ (.A(_04060_),
    .X(_00672_));
 sky130_fd_sc_hd__nand2_1 _19360_ (.A(_04042_),
    .B(_12238_),
    .Y(_04061_));
 sky130_fd_sc_hd__o211a_1 _19361_ (.A1(_03248_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__mux2_1 _19362_ (.A0(_04062_),
    .A1(net3781),
    .S(_04031_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _19363_ (.A(_04063_),
    .X(_00673_));
 sky130_fd_sc_hd__nand2_1 _19364_ (.A(_04042_),
    .B(_12246_),
    .Y(_04064_));
 sky130_fd_sc_hd__o211a_1 _19365_ (.A1(_03252_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__mux2_1 _19366_ (.A0(_04065_),
    .A1(net3630),
    .S(_04031_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _19367_ (.A(_04066_),
    .X(_00674_));
 sky130_fd_sc_hd__o211a_1 _19368_ (.A1(_03256_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04043_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_8 _19369_ (.A(_04030_),
    .X(_04068_));
 sky130_fd_sc_hd__mux2_1 _19370_ (.A0(_04067_),
    .A1(net3403),
    .S(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _19371_ (.A(_04069_),
    .X(_00675_));
 sky130_fd_sc_hd__o211a_1 _19372_ (.A1(_03261_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04046_),
    .X(_04070_));
 sky130_fd_sc_hd__mux2_1 _19373_ (.A0(_04070_),
    .A1(net2438),
    .S(_04068_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _19374_ (.A(_04071_),
    .X(_00676_));
 sky130_fd_sc_hd__o211a_1 _19375_ (.A1(_03264_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04049_),
    .X(_04072_));
 sky130_fd_sc_hd__mux2_1 _19376_ (.A0(_04072_),
    .A1(net3115),
    .S(_04068_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_1 _19377_ (.A(_04073_),
    .X(_00677_));
 sky130_fd_sc_hd__o211a_1 _19378_ (.A1(_03267_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04052_),
    .X(_04074_));
 sky130_fd_sc_hd__mux2_1 _19379_ (.A0(_04074_),
    .A1(net3040),
    .S(_04068_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _19380_ (.A(_04075_),
    .X(_00678_));
 sky130_fd_sc_hd__o211a_1 _19381_ (.A1(_03270_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04055_),
    .X(_04076_));
 sky130_fd_sc_hd__mux2_1 _19382_ (.A0(_04076_),
    .A1(net2734),
    .S(_04068_),
    .X(_04077_));
 sky130_fd_sc_hd__clkbuf_1 _19383_ (.A(_04077_),
    .X(_00679_));
 sky130_fd_sc_hd__o211a_1 _19384_ (.A1(_03273_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04058_),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_1 _19385_ (.A0(_04078_),
    .A1(net3581),
    .S(_04068_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _19386_ (.A(_04079_),
    .X(_00680_));
 sky130_fd_sc_hd__o211a_1 _19387_ (.A1(_03276_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04061_),
    .X(_04080_));
 sky130_fd_sc_hd__mux2_1 _19388_ (.A0(_04080_),
    .A1(net2389),
    .S(_04068_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _19389_ (.A(_04081_),
    .X(_00681_));
 sky130_fd_sc_hd__o211a_1 _19390_ (.A1(_03279_),
    .A2(_04040_),
    .B1(_04041_),
    .C1(_04064_),
    .X(_04082_));
 sky130_fd_sc_hd__mux2_1 _19391_ (.A0(_04082_),
    .A1(net2664),
    .S(_04068_),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _19392_ (.A(_04083_),
    .X(_00682_));
 sky130_fd_sc_hd__clkbuf_8 _19393_ (.A(_03702_),
    .X(_04084_));
 sky130_fd_sc_hd__o211a_1 _19394_ (.A1(_12170_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04043_),
    .X(_04085_));
 sky130_fd_sc_hd__mux2_1 _19395_ (.A0(_04085_),
    .A1(net2178),
    .S(_04068_),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _19396_ (.A(_04086_),
    .X(_00683_));
 sky130_fd_sc_hd__o211a_1 _19397_ (.A1(_12195_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04046_),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _19398_ (.A0(_04087_),
    .A1(net2081),
    .S(_04068_),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_1 _19399_ (.A(_04088_),
    .X(_00684_));
 sky130_fd_sc_hd__o211a_1 _19400_ (.A1(_12203_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04049_),
    .X(_04089_));
 sky130_fd_sc_hd__mux2_1 _19401_ (.A0(_04089_),
    .A1(net2046),
    .S(_04068_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _19402_ (.A(_04090_),
    .X(_00685_));
 sky130_fd_sc_hd__o211a_1 _19403_ (.A1(_12211_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04052_),
    .X(_04091_));
 sky130_fd_sc_hd__mux2_1 _19404_ (.A0(_04091_),
    .A1(net2036),
    .S(_04068_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _19405_ (.A(_04092_),
    .X(_00686_));
 sky130_fd_sc_hd__o211a_1 _19406_ (.A1(_12219_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04055_),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_1 _19407_ (.A0(_04093_),
    .A1(net2370),
    .S(_04068_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _19408_ (.A(_04094_),
    .X(_00687_));
 sky130_fd_sc_hd__o211a_1 _19409_ (.A1(_12227_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04058_),
    .X(_04095_));
 sky130_fd_sc_hd__mux2_1 _19410_ (.A0(_04095_),
    .A1(net2291),
    .S(_04068_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _19411_ (.A(_04096_),
    .X(_00688_));
 sky130_fd_sc_hd__o211a_1 _19412_ (.A1(_12235_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04061_),
    .X(_04097_));
 sky130_fd_sc_hd__mux2_1 _19413_ (.A0(_04097_),
    .A1(net2097),
    .S(_04068_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _19414_ (.A(_04098_),
    .X(_00689_));
 sky130_fd_sc_hd__o211a_1 _19415_ (.A1(_12243_),
    .A2(_04042_),
    .B1(_04084_),
    .C1(_04064_),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _19416_ (.A0(_04099_),
    .A1(net2059),
    .S(_04068_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _19417_ (.A(_04100_),
    .X(_00690_));
 sky130_fd_sc_hd__clkbuf_8 _19418_ (.A(_02809_),
    .X(_04101_));
 sky130_fd_sc_hd__inv_2 _19419_ (.A(\line_cache_idx[7] ),
    .Y(_04102_));
 sky130_fd_sc_hd__and3_4 _19420_ (.A(_02813_),
    .B(_04102_),
    .C(\line_cache_idx[6] ),
    .X(_04103_));
 sky130_fd_sc_hd__nor2_8 _19421_ (.A(_09070_),
    .B(_02812_),
    .Y(_04104_));
 sky130_fd_sc_hd__nand2_1 _19422_ (.A(_04103_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__a21bo_1 _19423_ (.A1(_04105_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_8 _19424_ (.A(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__mux2_1 _19425_ (.A0(_04101_),
    .A1(net2918),
    .S(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _19426_ (.A(_04108_),
    .X(_00691_));
 sky130_fd_sc_hd__buf_6 _19427_ (.A(_02822_),
    .X(_04109_));
 sky130_fd_sc_hd__mux2_1 _19428_ (.A0(_04109_),
    .A1(net2690),
    .S(_04107_),
    .X(_04110_));
 sky130_fd_sc_hd__clkbuf_1 _19429_ (.A(_04110_),
    .X(_00692_));
 sky130_fd_sc_hd__buf_8 _19430_ (.A(_02826_),
    .X(_04111_));
 sky130_fd_sc_hd__mux2_1 _19431_ (.A0(_04111_),
    .A1(net3415),
    .S(_04107_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _19432_ (.A(_04112_),
    .X(_00693_));
 sky130_fd_sc_hd__buf_8 _19433_ (.A(_02830_),
    .X(_04113_));
 sky130_fd_sc_hd__mux2_1 _19434_ (.A0(_04113_),
    .A1(net2545),
    .S(_04107_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _19435_ (.A(_04114_),
    .X(_00694_));
 sky130_fd_sc_hd__buf_8 _19436_ (.A(_02834_),
    .X(_04115_));
 sky130_fd_sc_hd__mux2_1 _19437_ (.A0(_04115_),
    .A1(net2989),
    .S(_04107_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _19438_ (.A(_04116_),
    .X(_00695_));
 sky130_fd_sc_hd__buf_8 _19439_ (.A(_02838_),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _19440_ (.A0(_04117_),
    .A1(net3357),
    .S(_04107_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _19441_ (.A(_04118_),
    .X(_00696_));
 sky130_fd_sc_hd__buf_8 _19442_ (.A(_02842_),
    .X(_04119_));
 sky130_fd_sc_hd__mux2_1 _19443_ (.A0(_04119_),
    .A1(net3246),
    .S(_04107_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _19444_ (.A(_04120_),
    .X(_00697_));
 sky130_fd_sc_hd__buf_8 _19445_ (.A(_02846_),
    .X(_04121_));
 sky130_fd_sc_hd__mux2_1 _19446_ (.A0(_04121_),
    .A1(net2530),
    .S(_04107_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _19447_ (.A(_04122_),
    .X(_00698_));
 sky130_fd_sc_hd__buf_4 _19448_ (.A(_04105_),
    .X(_04123_));
 sky130_fd_sc_hd__buf_4 _19449_ (.A(_04105_),
    .X(_04124_));
 sky130_fd_sc_hd__nand2_1 _19450_ (.A(_04124_),
    .B(_12185_),
    .Y(_04125_));
 sky130_fd_sc_hd__o211a_1 _19451_ (.A1(_03222_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__mux2_1 _19452_ (.A0(_04126_),
    .A1(net2319),
    .S(_04107_),
    .X(_04127_));
 sky130_fd_sc_hd__clkbuf_1 _19453_ (.A(_04127_),
    .X(_00699_));
 sky130_fd_sc_hd__nand2_1 _19454_ (.A(_04124_),
    .B(_12198_),
    .Y(_04128_));
 sky130_fd_sc_hd__o211a_1 _19455_ (.A1(_03228_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__mux2_1 _19456_ (.A0(_04129_),
    .A1(net2221),
    .S(_04107_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _19457_ (.A(_04130_),
    .X(_00700_));
 sky130_fd_sc_hd__nand2_1 _19458_ (.A(_04124_),
    .B(_12206_),
    .Y(_04131_));
 sky130_fd_sc_hd__o211a_1 _19459_ (.A1(_03232_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__mux2_1 _19460_ (.A0(_04132_),
    .A1(net2610),
    .S(_04107_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _19461_ (.A(_04133_),
    .X(_00701_));
 sky130_fd_sc_hd__nand2_1 _19462_ (.A(_04124_),
    .B(_12214_),
    .Y(_04134_));
 sky130_fd_sc_hd__o211a_1 _19463_ (.A1(_03236_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__mux2_1 _19464_ (.A0(_04135_),
    .A1(net2854),
    .S(_04107_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _19465_ (.A(_04136_),
    .X(_00702_));
 sky130_fd_sc_hd__nand2_1 _19466_ (.A(_04124_),
    .B(_12222_),
    .Y(_04137_));
 sky130_fd_sc_hd__o211a_1 _19467_ (.A1(_03240_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__mux2_1 _19468_ (.A0(_04138_),
    .A1(net2737),
    .S(_04107_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _19469_ (.A(_04139_),
    .X(_00703_));
 sky130_fd_sc_hd__nand2_1 _19470_ (.A(_04124_),
    .B(_12230_),
    .Y(_04140_));
 sky130_fd_sc_hd__o211a_1 _19471_ (.A1(_03244_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__mux2_1 _19472_ (.A0(_04141_),
    .A1(net3122),
    .S(_04107_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _19473_ (.A(_04142_),
    .X(_00704_));
 sky130_fd_sc_hd__nand2_1 _19474_ (.A(_04124_),
    .B(_12238_),
    .Y(_04143_));
 sky130_fd_sc_hd__o211a_1 _19475_ (.A1(_03248_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__mux2_1 _19476_ (.A0(_04144_),
    .A1(net2372),
    .S(_04107_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _19477_ (.A(_04145_),
    .X(_00705_));
 sky130_fd_sc_hd__nand2_1 _19478_ (.A(_04124_),
    .B(_12246_),
    .Y(_04146_));
 sky130_fd_sc_hd__o211a_1 _19479_ (.A1(_03252_),
    .A2(_04123_),
    .B1(_04084_),
    .C1(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__mux2_1 _19480_ (.A0(_04147_),
    .A1(net2870),
    .S(_04107_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_1 _19481_ (.A(_04148_),
    .X(_00706_));
 sky130_fd_sc_hd__buf_4 _19482_ (.A(_03702_),
    .X(_04149_));
 sky130_fd_sc_hd__o211a_1 _19483_ (.A1(_03256_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04125_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_8 _19484_ (.A(_04106_),
    .X(_04151_));
 sky130_fd_sc_hd__mux2_1 _19485_ (.A0(_04150_),
    .A1(net2725),
    .S(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _19486_ (.A(_04152_),
    .X(_00707_));
 sky130_fd_sc_hd__o211a_1 _19487_ (.A1(_03261_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04128_),
    .X(_04153_));
 sky130_fd_sc_hd__mux2_1 _19488_ (.A0(_04153_),
    .A1(net2656),
    .S(_04151_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _19489_ (.A(_04154_),
    .X(_00708_));
 sky130_fd_sc_hd__o211a_1 _19490_ (.A1(_03264_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04131_),
    .X(_04155_));
 sky130_fd_sc_hd__mux2_1 _19491_ (.A0(_04155_),
    .A1(net2905),
    .S(_04151_),
    .X(_04156_));
 sky130_fd_sc_hd__clkbuf_1 _19492_ (.A(_04156_),
    .X(_00709_));
 sky130_fd_sc_hd__o211a_1 _19493_ (.A1(_03267_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04134_),
    .X(_04157_));
 sky130_fd_sc_hd__mux2_1 _19494_ (.A0(_04157_),
    .A1(net3118),
    .S(_04151_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _19495_ (.A(_04158_),
    .X(_00710_));
 sky130_fd_sc_hd__o211a_1 _19496_ (.A1(_03270_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04137_),
    .X(_04159_));
 sky130_fd_sc_hd__mux2_1 _19497_ (.A0(_04159_),
    .A1(net3345),
    .S(_04151_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _19498_ (.A(_04160_),
    .X(_00711_));
 sky130_fd_sc_hd__o211a_1 _19499_ (.A1(_03273_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04140_),
    .X(_04161_));
 sky130_fd_sc_hd__mux2_1 _19500_ (.A0(_04161_),
    .A1(net2745),
    .S(_04151_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _19501_ (.A(_04162_),
    .X(_00712_));
 sky130_fd_sc_hd__o211a_1 _19502_ (.A1(_03276_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04143_),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_1 _19503_ (.A0(_04163_),
    .A1(net3221),
    .S(_04151_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _19504_ (.A(_04164_),
    .X(_00713_));
 sky130_fd_sc_hd__o211a_1 _19505_ (.A1(_03279_),
    .A2(_04123_),
    .B1(_04149_),
    .C1(_04146_),
    .X(_04165_));
 sky130_fd_sc_hd__mux2_1 _19506_ (.A0(_04165_),
    .A1(net2958),
    .S(_04151_),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _19507_ (.A(_04166_),
    .X(_00714_));
 sky130_fd_sc_hd__o211a_1 _19508_ (.A1(_12170_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04125_),
    .X(_04167_));
 sky130_fd_sc_hd__mux2_1 _19509_ (.A0(_04167_),
    .A1(net3008),
    .S(_04151_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _19510_ (.A(_04168_),
    .X(_00715_));
 sky130_fd_sc_hd__o211a_1 _19511_ (.A1(_12195_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04128_),
    .X(_04169_));
 sky130_fd_sc_hd__mux2_1 _19512_ (.A0(_04169_),
    .A1(net3090),
    .S(_04151_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_1 _19513_ (.A(_04170_),
    .X(_00716_));
 sky130_fd_sc_hd__o211a_1 _19514_ (.A1(_12203_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04131_),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _19515_ (.A0(_04171_),
    .A1(net3394),
    .S(_04151_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _19516_ (.A(_04172_),
    .X(_00717_));
 sky130_fd_sc_hd__o211a_1 _19517_ (.A1(_12211_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04134_),
    .X(_04173_));
 sky130_fd_sc_hd__mux2_1 _19518_ (.A0(_04173_),
    .A1(net3361),
    .S(_04151_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _19519_ (.A(_04174_),
    .X(_00718_));
 sky130_fd_sc_hd__o211a_1 _19520_ (.A1(_12219_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04137_),
    .X(_04175_));
 sky130_fd_sc_hd__mux2_1 _19521_ (.A0(_04175_),
    .A1(net3399),
    .S(_04151_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _19522_ (.A(_04176_),
    .X(_00719_));
 sky130_fd_sc_hd__o211a_1 _19523_ (.A1(_12227_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04140_),
    .X(_04177_));
 sky130_fd_sc_hd__mux2_1 _19524_ (.A0(_04177_),
    .A1(net3456),
    .S(_04151_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _19525_ (.A(_04178_),
    .X(_00720_));
 sky130_fd_sc_hd__o211a_1 _19526_ (.A1(_12235_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04143_),
    .X(_04179_));
 sky130_fd_sc_hd__mux2_1 _19527_ (.A0(_04179_),
    .A1(net3294),
    .S(_04151_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _19528_ (.A(_04180_),
    .X(_00721_));
 sky130_fd_sc_hd__o211a_1 _19529_ (.A1(_12243_),
    .A2(_04124_),
    .B1(_04149_),
    .C1(_04146_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _19530_ (.A0(_04181_),
    .A1(net2161),
    .S(_04151_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _19531_ (.A(_04182_),
    .X(_00722_));
 sky130_fd_sc_hd__nor2_8 _19532_ (.A(_09070_),
    .B(_12293_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _19533_ (.A(_04103_),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__inv_2 _19534_ (.A(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__o21ai_4 _19535_ (.A1(_12290_),
    .A2(_04185_),
    .B1(_02818_),
    .Y(_04186_));
 sky130_fd_sc_hd__mux2_1 _19536_ (.A0(_04101_),
    .A1(net2761),
    .S(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _19537_ (.A(_04187_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _19538_ (.A0(_04109_),
    .A1(net3396),
    .S(_04186_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _19539_ (.A(_04188_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _19540_ (.A0(_04111_),
    .A1(net3492),
    .S(_04186_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _19541_ (.A(_04189_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _19542_ (.A0(_04113_),
    .A1(net2290),
    .S(_04186_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _19543_ (.A(_04190_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _19544_ (.A0(_04115_),
    .A1(net3421),
    .S(_04186_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _19545_ (.A(_04191_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _19546_ (.A0(_04117_),
    .A1(net2495),
    .S(_04186_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _19547_ (.A(_04192_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _19548_ (.A0(_04119_),
    .A1(net2696),
    .S(_04186_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _19549_ (.A(_04193_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _19550_ (.A0(_04121_),
    .A1(net2600),
    .S(_04186_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _19551_ (.A(_04194_),
    .X(_00730_));
 sky130_fd_sc_hd__buf_4 _19552_ (.A(_04186_),
    .X(_04195_));
 sky130_fd_sc_hd__buf_4 _19553_ (.A(_04185_),
    .X(_04196_));
 sky130_fd_sc_hd__buf_4 _19554_ (.A(_04185_),
    .X(_04197_));
 sky130_fd_sc_hd__nor2_1 _19555_ (.A(_02854_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__a211o_1 _19556_ (.A1(_02852_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__buf_4 _19557_ (.A(_04186_),
    .X(_04200_));
 sky130_fd_sc_hd__nand2_1 _19558_ (.A(_04200_),
    .B(net976),
    .Y(_04201_));
 sky130_fd_sc_hd__o21ai_1 _19559_ (.A1(_04195_),
    .A2(_04199_),
    .B1(net977),
    .Y(_00731_));
 sky130_fd_sc_hd__nor2_1 _19560_ (.A(_02863_),
    .B(_04197_),
    .Y(_04202_));
 sky130_fd_sc_hd__a211o_1 _19561_ (.A1(_02862_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__nand2_1 _19562_ (.A(_04200_),
    .B(net508),
    .Y(_04204_));
 sky130_fd_sc_hd__o21ai_1 _19563_ (.A1(_04195_),
    .A2(_04203_),
    .B1(net509),
    .Y(_00732_));
 sky130_fd_sc_hd__nor2_1 _19564_ (.A(_02870_),
    .B(_04197_),
    .Y(_04205_));
 sky130_fd_sc_hd__a211o_1 _19565_ (.A1(_02869_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__nand2_1 _19566_ (.A(_04200_),
    .B(net1134),
    .Y(_04207_));
 sky130_fd_sc_hd__o21ai_1 _19567_ (.A1(_04195_),
    .A2(_04206_),
    .B1(net1135),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2_1 _19568_ (.A(_02877_),
    .B(_04197_),
    .Y(_04208_));
 sky130_fd_sc_hd__a211o_1 _19569_ (.A1(_02876_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__nand2_1 _19570_ (.A(_04200_),
    .B(net678),
    .Y(_04210_));
 sky130_fd_sc_hd__o21ai_1 _19571_ (.A1(_04195_),
    .A2(_04209_),
    .B1(net679),
    .Y(_00734_));
 sky130_fd_sc_hd__nor2_1 _19572_ (.A(_02884_),
    .B(_04197_),
    .Y(_04211_));
 sky130_fd_sc_hd__a211o_1 _19573_ (.A1(_02883_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__nand2_1 _19574_ (.A(_04200_),
    .B(net1100),
    .Y(_04213_));
 sky130_fd_sc_hd__o21ai_1 _19575_ (.A1(_04195_),
    .A2(_04212_),
    .B1(net1101),
    .Y(_00735_));
 sky130_fd_sc_hd__nor2_1 _19576_ (.A(_02891_),
    .B(_04197_),
    .Y(_04214_));
 sky130_fd_sc_hd__a211o_1 _19577_ (.A1(_02890_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__nand2_1 _19578_ (.A(_04200_),
    .B(net736),
    .Y(_04216_));
 sky130_fd_sc_hd__o21ai_1 _19579_ (.A1(_04195_),
    .A2(_04215_),
    .B1(net737),
    .Y(_00736_));
 sky130_fd_sc_hd__nor2_1 _19580_ (.A(_02898_),
    .B(_04197_),
    .Y(_04217_));
 sky130_fd_sc_hd__a211o_1 _19581_ (.A1(_02897_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__nand2_1 _19582_ (.A(_04200_),
    .B(net872),
    .Y(_04219_));
 sky130_fd_sc_hd__o21ai_1 _19583_ (.A1(_04195_),
    .A2(_04218_),
    .B1(net873),
    .Y(_00737_));
 sky130_fd_sc_hd__nor2_1 _19584_ (.A(_02905_),
    .B(_04197_),
    .Y(_04220_));
 sky130_fd_sc_hd__a211o_1 _19585_ (.A1(_02904_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__nand2_1 _19586_ (.A(_04200_),
    .B(net784),
    .Y(_04222_));
 sky130_fd_sc_hd__o21ai_1 _19587_ (.A1(_04195_),
    .A2(_04221_),
    .B1(net785),
    .Y(_00738_));
 sky130_fd_sc_hd__buf_4 _19588_ (.A(_04186_),
    .X(_04223_));
 sky130_fd_sc_hd__a211o_1 _19589_ (.A1(_02912_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04198_),
    .X(_04224_));
 sky130_fd_sc_hd__nand2_1 _19590_ (.A(_04200_),
    .B(net1422),
    .Y(_04225_));
 sky130_fd_sc_hd__o21ai_1 _19591_ (.A1(_04223_),
    .A2(_04224_),
    .B1(net1423),
    .Y(_00739_));
 sky130_fd_sc_hd__a211o_1 _19592_ (.A1(_02917_),
    .A2(_04196_),
    .B1(_03194_),
    .C1(_04202_),
    .X(_04226_));
 sky130_fd_sc_hd__nand2_1 _19593_ (.A(_04200_),
    .B(net604),
    .Y(_04227_));
 sky130_fd_sc_hd__o21ai_1 _19594_ (.A1(_04223_),
    .A2(_04226_),
    .B1(net605),
    .Y(_00740_));
 sky130_fd_sc_hd__buf_4 _19595_ (.A(_09129_),
    .X(_04228_));
 sky130_fd_sc_hd__a211o_1 _19596_ (.A1(_02922_),
    .A2(_04196_),
    .B1(_04228_),
    .C1(_04205_),
    .X(_04229_));
 sky130_fd_sc_hd__nand2_1 _19597_ (.A(_04200_),
    .B(net560),
    .Y(_04230_));
 sky130_fd_sc_hd__o21ai_1 _19598_ (.A1(_04223_),
    .A2(_04229_),
    .B1(net561),
    .Y(_00741_));
 sky130_fd_sc_hd__a211o_1 _19599_ (.A1(_02928_),
    .A2(_04196_),
    .B1(_04228_),
    .C1(_04208_),
    .X(_04231_));
 sky130_fd_sc_hd__nand2_1 _19600_ (.A(_04200_),
    .B(net468),
    .Y(_04232_));
 sky130_fd_sc_hd__o21ai_1 _19601_ (.A1(_04223_),
    .A2(_04231_),
    .B1(net469),
    .Y(_00742_));
 sky130_fd_sc_hd__a211o_1 _19602_ (.A1(_02933_),
    .A2(_04196_),
    .B1(_04228_),
    .C1(_04211_),
    .X(_04233_));
 sky130_fd_sc_hd__nand2_1 _19603_ (.A(_04200_),
    .B(net1206),
    .Y(_04234_));
 sky130_fd_sc_hd__o21ai_1 _19604_ (.A1(_04223_),
    .A2(_04233_),
    .B1(net1207),
    .Y(_00743_));
 sky130_fd_sc_hd__a211o_1 _19605_ (.A1(_02938_),
    .A2(_04196_),
    .B1(_04228_),
    .C1(_04214_),
    .X(_04235_));
 sky130_fd_sc_hd__nand2_1 _19606_ (.A(_04200_),
    .B(net822),
    .Y(_04236_));
 sky130_fd_sc_hd__o21ai_1 _19607_ (.A1(_04223_),
    .A2(_04235_),
    .B1(net823),
    .Y(_00744_));
 sky130_fd_sc_hd__a211o_1 _19608_ (.A1(_02943_),
    .A2(_04196_),
    .B1(_04228_),
    .C1(_04217_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _19609_ (.A(_04200_),
    .B(net1128),
    .Y(_04238_));
 sky130_fd_sc_hd__o21ai_1 _19610_ (.A1(_04223_),
    .A2(_04237_),
    .B1(net1129),
    .Y(_00745_));
 sky130_fd_sc_hd__a211o_1 _19611_ (.A1(_02948_),
    .A2(_04196_),
    .B1(_04228_),
    .C1(_04220_),
    .X(_04239_));
 sky130_fd_sc_hd__nand2_1 _19612_ (.A(_04200_),
    .B(net850),
    .Y(_04240_));
 sky130_fd_sc_hd__o21ai_1 _19613_ (.A1(_04223_),
    .A2(_04239_),
    .B1(net851),
    .Y(_00746_));
 sky130_fd_sc_hd__a211o_1 _19614_ (.A1(_02952_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04198_),
    .X(_04241_));
 sky130_fd_sc_hd__nand2_1 _19615_ (.A(_04195_),
    .B(net1286),
    .Y(_04242_));
 sky130_fd_sc_hd__o21ai_1 _19616_ (.A1(_04223_),
    .A2(_04241_),
    .B1(net1287),
    .Y(_00747_));
 sky130_fd_sc_hd__a211o_1 _19617_ (.A1(_02956_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04202_),
    .X(_04243_));
 sky130_fd_sc_hd__nand2_1 _19618_ (.A(_04195_),
    .B(net1626),
    .Y(_04244_));
 sky130_fd_sc_hd__o21ai_1 _19619_ (.A1(_04223_),
    .A2(_04243_),
    .B1(net1627),
    .Y(_00748_));
 sky130_fd_sc_hd__a211o_1 _19620_ (.A1(_02960_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04205_),
    .X(_04245_));
 sky130_fd_sc_hd__nand2_1 _19621_ (.A(_04195_),
    .B(net950),
    .Y(_04246_));
 sky130_fd_sc_hd__o21ai_1 _19622_ (.A1(_04223_),
    .A2(_04245_),
    .B1(net951),
    .Y(_00749_));
 sky130_fd_sc_hd__a211o_1 _19623_ (.A1(_02964_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04208_),
    .X(_04247_));
 sky130_fd_sc_hd__nand2_1 _19624_ (.A(_04195_),
    .B(net1814),
    .Y(_04248_));
 sky130_fd_sc_hd__o21ai_1 _19625_ (.A1(_04223_),
    .A2(_04247_),
    .B1(net1815),
    .Y(_00750_));
 sky130_fd_sc_hd__a211o_1 _19626_ (.A1(_02968_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04211_),
    .X(_04249_));
 sky130_fd_sc_hd__nand2_1 _19627_ (.A(_04195_),
    .B(net1736),
    .Y(_04250_));
 sky130_fd_sc_hd__o21ai_1 _19628_ (.A1(_04223_),
    .A2(_04249_),
    .B1(net1737),
    .Y(_00751_));
 sky130_fd_sc_hd__a211o_1 _19629_ (.A1(_02972_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04214_),
    .X(_04251_));
 sky130_fd_sc_hd__nand2_1 _19630_ (.A(_04195_),
    .B(net1885),
    .Y(_04252_));
 sky130_fd_sc_hd__o21ai_1 _19631_ (.A1(_04223_),
    .A2(_04251_),
    .B1(net1886),
    .Y(_00752_));
 sky130_fd_sc_hd__a211o_1 _19632_ (.A1(_02976_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04217_),
    .X(_04253_));
 sky130_fd_sc_hd__nand2_1 _19633_ (.A(_04195_),
    .B(net1792),
    .Y(_04254_));
 sky130_fd_sc_hd__o21ai_1 _19634_ (.A1(_04223_),
    .A2(_04253_),
    .B1(net1793),
    .Y(_00753_));
 sky130_fd_sc_hd__a211o_1 _19635_ (.A1(_02980_),
    .A2(_04197_),
    .B1(_04228_),
    .C1(_04220_),
    .X(_04255_));
 sky130_fd_sc_hd__nand2_1 _19636_ (.A(_04195_),
    .B(net1812),
    .Y(_04256_));
 sky130_fd_sc_hd__o21ai_1 _19637_ (.A1(_04223_),
    .A2(_04255_),
    .B1(net1813),
    .Y(_00754_));
 sky130_fd_sc_hd__nor2_8 _19638_ (.A(_09070_),
    .B(_12292_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_1 _19639_ (.A(_04103_),
    .B(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__inv_2 _19640_ (.A(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__o21ai_4 _19641_ (.A1(_12290_),
    .A2(_04259_),
    .B1(_02818_),
    .Y(_04260_));
 sky130_fd_sc_hd__mux2_1 _19642_ (.A0(_04101_),
    .A1(net3555),
    .S(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _19643_ (.A(_04261_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _19644_ (.A0(_04109_),
    .A1(net2489),
    .S(_04260_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _19645_ (.A(_04262_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _19646_ (.A0(_04111_),
    .A1(net3442),
    .S(_04260_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _19647_ (.A(_04263_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _19648_ (.A0(_04113_),
    .A1(net2535),
    .S(_04260_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _19649_ (.A(_04264_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _19650_ (.A0(_04115_),
    .A1(net3613),
    .S(_04260_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _19651_ (.A(_04265_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _19652_ (.A0(_04117_),
    .A1(net2238),
    .S(_04260_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _19653_ (.A(_04266_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _19654_ (.A0(_04119_),
    .A1(net3347),
    .S(_04260_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _19655_ (.A(_04267_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _19656_ (.A0(_04121_),
    .A1(net2727),
    .S(_04260_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _19657_ (.A(_04268_),
    .X(_00762_));
 sky130_fd_sc_hd__buf_4 _19658_ (.A(_04260_),
    .X(_04269_));
 sky130_fd_sc_hd__buf_4 _19659_ (.A(_04259_),
    .X(_04270_));
 sky130_fd_sc_hd__buf_4 _19660_ (.A(_04259_),
    .X(_04271_));
 sky130_fd_sc_hd__nor2_1 _19661_ (.A(_02854_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__a211o_1 _19662_ (.A1(_02852_),
    .A2(_04270_),
    .B1(_04228_),
    .C1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__buf_4 _19663_ (.A(_04260_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2_1 _19664_ (.A(_04274_),
    .B(net500),
    .Y(_04275_));
 sky130_fd_sc_hd__o21ai_1 _19665_ (.A1(_04269_),
    .A2(_04273_),
    .B1(net501),
    .Y(_00763_));
 sky130_fd_sc_hd__nor2_1 _19666_ (.A(_02863_),
    .B(_04271_),
    .Y(_04276_));
 sky130_fd_sc_hd__a211o_1 _19667_ (.A1(_02862_),
    .A2(_04270_),
    .B1(_04228_),
    .C1(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__nand2_1 _19668_ (.A(_04274_),
    .B(net486),
    .Y(_04278_));
 sky130_fd_sc_hd__o21ai_1 _19669_ (.A1(_04269_),
    .A2(_04277_),
    .B1(net487),
    .Y(_00764_));
 sky130_fd_sc_hd__buf_4 _19670_ (.A(_09129_),
    .X(_04279_));
 sky130_fd_sc_hd__nor2_1 _19671_ (.A(_02870_),
    .B(_04271_),
    .Y(_04280_));
 sky130_fd_sc_hd__a211o_1 _19672_ (.A1(_02869_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__nand2_1 _19673_ (.A(_04274_),
    .B(net480),
    .Y(_04282_));
 sky130_fd_sc_hd__o21ai_1 _19674_ (.A1(_04269_),
    .A2(_04281_),
    .B1(net481),
    .Y(_00765_));
 sky130_fd_sc_hd__nor2_1 _19675_ (.A(_02877_),
    .B(_04271_),
    .Y(_04283_));
 sky130_fd_sc_hd__a211o_1 _19676_ (.A1(_02876_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__nand2_1 _19677_ (.A(_04274_),
    .B(net518),
    .Y(_04285_));
 sky130_fd_sc_hd__o21ai_1 _19678_ (.A1(_04269_),
    .A2(_04284_),
    .B1(net519),
    .Y(_00766_));
 sky130_fd_sc_hd__nor2_1 _19679_ (.A(_02884_),
    .B(_04271_),
    .Y(_04286_));
 sky130_fd_sc_hd__a211o_1 _19680_ (.A1(_02883_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_1 _19681_ (.A(_04274_),
    .B(net1490),
    .Y(_04288_));
 sky130_fd_sc_hd__o21ai_1 _19682_ (.A1(_04269_),
    .A2(_04287_),
    .B1(net1491),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2_1 _19683_ (.A(_02891_),
    .B(_04271_),
    .Y(_04289_));
 sky130_fd_sc_hd__a211o_1 _19684_ (.A1(_02890_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04289_),
    .X(_04290_));
 sky130_fd_sc_hd__nand2_1 _19685_ (.A(_04274_),
    .B(net482),
    .Y(_04291_));
 sky130_fd_sc_hd__o21ai_1 _19686_ (.A1(_04269_),
    .A2(_04290_),
    .B1(net483),
    .Y(_00768_));
 sky130_fd_sc_hd__nor2_1 _19687_ (.A(_02898_),
    .B(_04271_),
    .Y(_04292_));
 sky130_fd_sc_hd__a211o_1 _19688_ (.A1(_02897_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__nand2_1 _19689_ (.A(_04274_),
    .B(net638),
    .Y(_04294_));
 sky130_fd_sc_hd__o21ai_1 _19690_ (.A1(_04269_),
    .A2(_04293_),
    .B1(net639),
    .Y(_00769_));
 sky130_fd_sc_hd__nor2_1 _19691_ (.A(_02905_),
    .B(_04271_),
    .Y(_04295_));
 sky130_fd_sc_hd__a211o_1 _19692_ (.A1(_02904_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__nand2_1 _19693_ (.A(_04274_),
    .B(net1324),
    .Y(_04297_));
 sky130_fd_sc_hd__o21ai_1 _19694_ (.A1(_04269_),
    .A2(_04296_),
    .B1(net1325),
    .Y(_00770_));
 sky130_fd_sc_hd__buf_4 _19695_ (.A(_04260_),
    .X(_04298_));
 sky130_fd_sc_hd__a211o_1 _19696_ (.A1(_02912_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04272_),
    .X(_04299_));
 sky130_fd_sc_hd__nand2_1 _19697_ (.A(_04274_),
    .B(net1226),
    .Y(_04300_));
 sky130_fd_sc_hd__o21ai_1 _19698_ (.A1(_04298_),
    .A2(_04299_),
    .B1(net1227),
    .Y(_00771_));
 sky130_fd_sc_hd__a211o_1 _19699_ (.A1(_02917_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04276_),
    .X(_04301_));
 sky130_fd_sc_hd__nand2_1 _19700_ (.A(_04274_),
    .B(net1500),
    .Y(_04302_));
 sky130_fd_sc_hd__o21ai_1 _19701_ (.A1(_04298_),
    .A2(_04301_),
    .B1(net1501),
    .Y(_00772_));
 sky130_fd_sc_hd__a211o_1 _19702_ (.A1(_02922_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04280_),
    .X(_04303_));
 sky130_fd_sc_hd__nand2_1 _19703_ (.A(_04274_),
    .B(net1842),
    .Y(_04304_));
 sky130_fd_sc_hd__o21ai_1 _19704_ (.A1(_04298_),
    .A2(_04303_),
    .B1(net1843),
    .Y(_00773_));
 sky130_fd_sc_hd__a211o_1 _19705_ (.A1(_02928_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04283_),
    .X(_04305_));
 sky130_fd_sc_hd__nand2_1 _19706_ (.A(_04274_),
    .B(net1716),
    .Y(_04306_));
 sky130_fd_sc_hd__o21ai_1 _19707_ (.A1(_04298_),
    .A2(_04305_),
    .B1(net1717),
    .Y(_00774_));
 sky130_fd_sc_hd__a211o_1 _19708_ (.A1(_02933_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04286_),
    .X(_04307_));
 sky130_fd_sc_hd__nand2_1 _19709_ (.A(_04274_),
    .B(net1688),
    .Y(_04308_));
 sky130_fd_sc_hd__o21ai_1 _19710_ (.A1(_04298_),
    .A2(_04307_),
    .B1(net1689),
    .Y(_00775_));
 sky130_fd_sc_hd__a211o_1 _19711_ (.A1(_02938_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04289_),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _19712_ (.A(_04274_),
    .B(net1534),
    .Y(_04310_));
 sky130_fd_sc_hd__o21ai_1 _19713_ (.A1(_04298_),
    .A2(_04309_),
    .B1(net1535),
    .Y(_00776_));
 sky130_fd_sc_hd__a211o_1 _19714_ (.A1(_02943_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04292_),
    .X(_04311_));
 sky130_fd_sc_hd__nand2_1 _19715_ (.A(_04274_),
    .B(net636),
    .Y(_04312_));
 sky130_fd_sc_hd__o21ai_1 _19716_ (.A1(_04298_),
    .A2(_04311_),
    .B1(net637),
    .Y(_00777_));
 sky130_fd_sc_hd__a211o_1 _19717_ (.A1(_02948_),
    .A2(_04270_),
    .B1(_04279_),
    .C1(_04295_),
    .X(_04313_));
 sky130_fd_sc_hd__nand2_1 _19718_ (.A(_04274_),
    .B(net916),
    .Y(_04314_));
 sky130_fd_sc_hd__o21ai_1 _19719_ (.A1(_04298_),
    .A2(_04313_),
    .B1(net917),
    .Y(_00778_));
 sky130_fd_sc_hd__a211o_1 _19720_ (.A1(_02952_),
    .A2(_04271_),
    .B1(_04279_),
    .C1(_04272_),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _19721_ (.A(_04269_),
    .B(net1760),
    .Y(_04316_));
 sky130_fd_sc_hd__o21ai_1 _19722_ (.A1(_04298_),
    .A2(_04315_),
    .B1(net1761),
    .Y(_00779_));
 sky130_fd_sc_hd__a211o_1 _19723_ (.A1(_02956_),
    .A2(_04271_),
    .B1(_04279_),
    .C1(_04276_),
    .X(_04317_));
 sky130_fd_sc_hd__nand2_1 _19724_ (.A(_04269_),
    .B(net1702),
    .Y(_04318_));
 sky130_fd_sc_hd__o21ai_1 _19725_ (.A1(_04298_),
    .A2(_04317_),
    .B1(net1703),
    .Y(_00780_));
 sky130_fd_sc_hd__buf_4 _19726_ (.A(_09129_),
    .X(_04319_));
 sky130_fd_sc_hd__a211o_1 _19727_ (.A1(_02960_),
    .A2(_04271_),
    .B1(_04319_),
    .C1(_04280_),
    .X(_04320_));
 sky130_fd_sc_hd__nand2_1 _19728_ (.A(_04269_),
    .B(net1822),
    .Y(_04321_));
 sky130_fd_sc_hd__o21ai_1 _19729_ (.A1(_04298_),
    .A2(_04320_),
    .B1(net1823),
    .Y(_00781_));
 sky130_fd_sc_hd__a211o_1 _19730_ (.A1(_02964_),
    .A2(_04271_),
    .B1(_04319_),
    .C1(_04283_),
    .X(_04322_));
 sky130_fd_sc_hd__nand2_1 _19731_ (.A(_04269_),
    .B(net1746),
    .Y(_04323_));
 sky130_fd_sc_hd__o21ai_1 _19732_ (.A1(_04298_),
    .A2(_04322_),
    .B1(net1747),
    .Y(_00782_));
 sky130_fd_sc_hd__a211o_1 _19733_ (.A1(_02968_),
    .A2(_04271_),
    .B1(_04319_),
    .C1(_04286_),
    .X(_04324_));
 sky130_fd_sc_hd__nand2_1 _19734_ (.A(_04269_),
    .B(net798),
    .Y(_04325_));
 sky130_fd_sc_hd__o21ai_1 _19735_ (.A1(_04298_),
    .A2(_04324_),
    .B1(net799),
    .Y(_00783_));
 sky130_fd_sc_hd__a211o_1 _19736_ (.A1(_02972_),
    .A2(_04271_),
    .B1(_04319_),
    .C1(_04289_),
    .X(_04326_));
 sky130_fd_sc_hd__nand2_1 _19737_ (.A(_04269_),
    .B(net1034),
    .Y(_04327_));
 sky130_fd_sc_hd__o21ai_1 _19738_ (.A1(_04298_),
    .A2(_04326_),
    .B1(net1035),
    .Y(_00784_));
 sky130_fd_sc_hd__a211o_1 _19739_ (.A1(_02976_),
    .A2(_04271_),
    .B1(_04319_),
    .C1(_04292_),
    .X(_04328_));
 sky130_fd_sc_hd__nand2_1 _19740_ (.A(_04269_),
    .B(net888),
    .Y(_04329_));
 sky130_fd_sc_hd__o21ai_1 _19741_ (.A1(_04298_),
    .A2(_04328_),
    .B1(net889),
    .Y(_00785_));
 sky130_fd_sc_hd__a211o_1 _19742_ (.A1(_02980_),
    .A2(_04271_),
    .B1(_04319_),
    .C1(_04295_),
    .X(_04330_));
 sky130_fd_sc_hd__nand2_1 _19743_ (.A(_04269_),
    .B(net724),
    .Y(_04331_));
 sky130_fd_sc_hd__o21ai_1 _19744_ (.A1(_04298_),
    .A2(_04330_),
    .B1(net725),
    .Y(_00786_));
 sky130_fd_sc_hd__clkbuf_16 _19745_ (.A(_12289_),
    .X(_04332_));
 sky130_fd_sc_hd__nor2_8 _19746_ (.A(_09070_),
    .B(_12171_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand2_1 _19747_ (.A(_04103_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__inv_2 _19748_ (.A(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__o21ai_4 _19749_ (.A1(_04332_),
    .A2(_04335_),
    .B1(_02818_),
    .Y(_04336_));
 sky130_fd_sc_hd__mux2_1 _19750_ (.A0(_04101_),
    .A1(net2056),
    .S(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _19751_ (.A(_04337_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _19752_ (.A0(_04109_),
    .A1(net2037),
    .S(_04336_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _19753_ (.A(_04338_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _19754_ (.A0(_04111_),
    .A1(net2086),
    .S(_04336_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _19755_ (.A(_04339_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _19756_ (.A0(_04113_),
    .A1(net2051),
    .S(_04336_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _19757_ (.A(_04340_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _19758_ (.A0(_04115_),
    .A1(net3406),
    .S(_04336_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _19759_ (.A(_04341_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _19760_ (.A0(_04117_),
    .A1(net2753),
    .S(_04336_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _19761_ (.A(_04342_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _19762_ (.A0(_04119_),
    .A1(net2126),
    .S(_04336_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _19763_ (.A(_04343_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _19764_ (.A0(_04121_),
    .A1(net2218),
    .S(_04336_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _19765_ (.A(_04344_),
    .X(_00794_));
 sky130_fd_sc_hd__buf_4 _19766_ (.A(_04336_),
    .X(_04345_));
 sky130_fd_sc_hd__buf_4 _19767_ (.A(_04335_),
    .X(_04346_));
 sky130_fd_sc_hd__buf_4 _19768_ (.A(_04335_),
    .X(_04347_));
 sky130_fd_sc_hd__nor2_1 _19769_ (.A(_02854_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__a211o_1 _19770_ (.A1(_02852_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__buf_4 _19771_ (.A(_04336_),
    .X(_04350_));
 sky130_fd_sc_hd__nand2_1 _19772_ (.A(_04350_),
    .B(net514),
    .Y(_04351_));
 sky130_fd_sc_hd__o21ai_1 _19773_ (.A1(_04345_),
    .A2(_04349_),
    .B1(net515),
    .Y(_00795_));
 sky130_fd_sc_hd__nor2_1 _19774_ (.A(_02863_),
    .B(_04347_),
    .Y(_04352_));
 sky130_fd_sc_hd__a211o_1 _19775_ (.A1(_02862_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__nand2_1 _19776_ (.A(_04350_),
    .B(net516),
    .Y(_04354_));
 sky130_fd_sc_hd__o21ai_1 _19777_ (.A1(_04345_),
    .A2(_04353_),
    .B1(net517),
    .Y(_00796_));
 sky130_fd_sc_hd__nor2_1 _19778_ (.A(_02870_),
    .B(_04347_),
    .Y(_04355_));
 sky130_fd_sc_hd__a211o_1 _19779_ (.A1(_02869_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__nand2_1 _19780_ (.A(_04350_),
    .B(net908),
    .Y(_04357_));
 sky130_fd_sc_hd__o21ai_1 _19781_ (.A1(_04345_),
    .A2(_04356_),
    .B1(net909),
    .Y(_00797_));
 sky130_fd_sc_hd__nor2_1 _19782_ (.A(_02877_),
    .B(_04347_),
    .Y(_04358_));
 sky130_fd_sc_hd__a211o_1 _19783_ (.A1(_02876_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__nand2_1 _19784_ (.A(_04350_),
    .B(net1150),
    .Y(_04360_));
 sky130_fd_sc_hd__o21ai_1 _19785_ (.A1(_04345_),
    .A2(_04359_),
    .B1(net1151),
    .Y(_00798_));
 sky130_fd_sc_hd__nor2_1 _19786_ (.A(_02884_),
    .B(_04347_),
    .Y(_04361_));
 sky130_fd_sc_hd__a211o_1 _19787_ (.A1(_02883_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__nand2_1 _19788_ (.A(_04350_),
    .B(net434),
    .Y(_04363_));
 sky130_fd_sc_hd__o21ai_1 _19789_ (.A1(_04345_),
    .A2(_04362_),
    .B1(net435),
    .Y(_00799_));
 sky130_fd_sc_hd__nor2_1 _19790_ (.A(_02891_),
    .B(_04347_),
    .Y(_04364_));
 sky130_fd_sc_hd__a211o_1 _19791_ (.A1(_02890_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__nand2_1 _19792_ (.A(_04350_),
    .B(net1740),
    .Y(_04366_));
 sky130_fd_sc_hd__o21ai_1 _19793_ (.A1(_04345_),
    .A2(_04365_),
    .B1(net1741),
    .Y(_00800_));
 sky130_fd_sc_hd__nor2_1 _19794_ (.A(_02898_),
    .B(_04347_),
    .Y(_04367_));
 sky130_fd_sc_hd__a211o_1 _19795_ (.A1(_02897_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__nand2_1 _19796_ (.A(_04350_),
    .B(net540),
    .Y(_04369_));
 sky130_fd_sc_hd__o21ai_1 _19797_ (.A1(_04345_),
    .A2(_04368_),
    .B1(net541),
    .Y(_00801_));
 sky130_fd_sc_hd__nor2_1 _19798_ (.A(_02905_),
    .B(_04347_),
    .Y(_04370_));
 sky130_fd_sc_hd__a211o_1 _19799_ (.A1(_02904_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__nand2_1 _19800_ (.A(_04350_),
    .B(net402),
    .Y(_04372_));
 sky130_fd_sc_hd__o21ai_1 _19801_ (.A1(_04345_),
    .A2(_04371_),
    .B1(net403),
    .Y(_00802_));
 sky130_fd_sc_hd__buf_4 _19802_ (.A(_04336_),
    .X(_04373_));
 sky130_fd_sc_hd__a211o_1 _19803_ (.A1(_02912_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04348_),
    .X(_04374_));
 sky130_fd_sc_hd__nand2_1 _19804_ (.A(_04350_),
    .B(net998),
    .Y(_04375_));
 sky130_fd_sc_hd__o21ai_1 _19805_ (.A1(_04373_),
    .A2(_04374_),
    .B1(net999),
    .Y(_00803_));
 sky130_fd_sc_hd__a211o_1 _19806_ (.A1(_02917_),
    .A2(_04346_),
    .B1(_04319_),
    .C1(_04352_),
    .X(_04376_));
 sky130_fd_sc_hd__nand2_1 _19807_ (.A(_04350_),
    .B(net474),
    .Y(_04377_));
 sky130_fd_sc_hd__o21ai_1 _19808_ (.A1(_04373_),
    .A2(_04376_),
    .B1(net475),
    .Y(_00804_));
 sky130_fd_sc_hd__buf_4 _19809_ (.A(_09129_),
    .X(_04378_));
 sky130_fd_sc_hd__a211o_1 _19810_ (.A1(_02922_),
    .A2(_04346_),
    .B1(_04378_),
    .C1(_04355_),
    .X(_04379_));
 sky130_fd_sc_hd__nand2_1 _19811_ (.A(_04350_),
    .B(net410),
    .Y(_04380_));
 sky130_fd_sc_hd__o21ai_1 _19812_ (.A1(_04373_),
    .A2(_04379_),
    .B1(net411),
    .Y(_00805_));
 sky130_fd_sc_hd__a211o_1 _19813_ (.A1(_02928_),
    .A2(_04346_),
    .B1(_04378_),
    .C1(_04358_),
    .X(_04381_));
 sky130_fd_sc_hd__nand2_1 _19814_ (.A(_04350_),
    .B(net408),
    .Y(_04382_));
 sky130_fd_sc_hd__o21ai_1 _19815_ (.A1(_04373_),
    .A2(_04381_),
    .B1(net409),
    .Y(_00806_));
 sky130_fd_sc_hd__a211o_1 _19816_ (.A1(_02933_),
    .A2(_04346_),
    .B1(_04378_),
    .C1(_04361_),
    .X(_04383_));
 sky130_fd_sc_hd__nand2_1 _19817_ (.A(_04350_),
    .B(net412),
    .Y(_04384_));
 sky130_fd_sc_hd__o21ai_1 _19818_ (.A1(_04373_),
    .A2(_04383_),
    .B1(net413),
    .Y(_00807_));
 sky130_fd_sc_hd__a211o_1 _19819_ (.A1(_02938_),
    .A2(_04346_),
    .B1(_04378_),
    .C1(_04364_),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_1 _19820_ (.A(_04350_),
    .B(net968),
    .Y(_04386_));
 sky130_fd_sc_hd__o21ai_1 _19821_ (.A1(_04373_),
    .A2(_04385_),
    .B1(net969),
    .Y(_00808_));
 sky130_fd_sc_hd__a211o_1 _19822_ (.A1(_02943_),
    .A2(_04346_),
    .B1(_04378_),
    .C1(_04367_),
    .X(_04387_));
 sky130_fd_sc_hd__nand2_1 _19823_ (.A(_04350_),
    .B(net396),
    .Y(_04388_));
 sky130_fd_sc_hd__o21ai_1 _19824_ (.A1(_04373_),
    .A2(_04387_),
    .B1(net397),
    .Y(_00809_));
 sky130_fd_sc_hd__a211o_1 _19825_ (.A1(_02948_),
    .A2(_04346_),
    .B1(_04378_),
    .C1(_04370_),
    .X(_04389_));
 sky130_fd_sc_hd__nand2_1 _19826_ (.A(_04350_),
    .B(net400),
    .Y(_04390_));
 sky130_fd_sc_hd__o21ai_1 _19827_ (.A1(_04373_),
    .A2(_04389_),
    .B1(net401),
    .Y(_00810_));
 sky130_fd_sc_hd__a211o_1 _19828_ (.A1(_02952_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04348_),
    .X(_04391_));
 sky130_fd_sc_hd__nand2_1 _19829_ (.A(_04345_),
    .B(net946),
    .Y(_04392_));
 sky130_fd_sc_hd__o21ai_1 _19830_ (.A1(_04373_),
    .A2(_04391_),
    .B1(net947),
    .Y(_00811_));
 sky130_fd_sc_hd__a211o_1 _19831_ (.A1(_02956_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04352_),
    .X(_04393_));
 sky130_fd_sc_hd__nand2_1 _19832_ (.A(_04345_),
    .B(net1524),
    .Y(_04394_));
 sky130_fd_sc_hd__o21ai_1 _19833_ (.A1(_04373_),
    .A2(_04393_),
    .B1(net1525),
    .Y(_00812_));
 sky130_fd_sc_hd__a211o_1 _19834_ (.A1(_02960_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04355_),
    .X(_04395_));
 sky130_fd_sc_hd__nand2_1 _19835_ (.A(_04345_),
    .B(net1348),
    .Y(_04396_));
 sky130_fd_sc_hd__o21ai_1 _19836_ (.A1(_04373_),
    .A2(_04395_),
    .B1(net1349),
    .Y(_00813_));
 sky130_fd_sc_hd__a211o_1 _19837_ (.A1(_02964_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04358_),
    .X(_04397_));
 sky130_fd_sc_hd__nand2_1 _19838_ (.A(_04345_),
    .B(net1336),
    .Y(_04398_));
 sky130_fd_sc_hd__o21ai_1 _19839_ (.A1(_04373_),
    .A2(_04397_),
    .B1(net1337),
    .Y(_00814_));
 sky130_fd_sc_hd__a211o_1 _19840_ (.A1(_02968_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04361_),
    .X(_04399_));
 sky130_fd_sc_hd__nand2_1 _19841_ (.A(_04345_),
    .B(net1212),
    .Y(_04400_));
 sky130_fd_sc_hd__o21ai_1 _19842_ (.A1(_04373_),
    .A2(_04399_),
    .B1(net1213),
    .Y(_00815_));
 sky130_fd_sc_hd__a211o_1 _19843_ (.A1(_02972_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04364_),
    .X(_04401_));
 sky130_fd_sc_hd__nand2_1 _19844_ (.A(_04345_),
    .B(net1272),
    .Y(_04402_));
 sky130_fd_sc_hd__o21ai_1 _19845_ (.A1(_04373_),
    .A2(_04401_),
    .B1(net1273),
    .Y(_00816_));
 sky130_fd_sc_hd__a211o_1 _19846_ (.A1(_02976_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04367_),
    .X(_04403_));
 sky130_fd_sc_hd__nand2_1 _19847_ (.A(_04345_),
    .B(net1552),
    .Y(_04404_));
 sky130_fd_sc_hd__o21ai_1 _19848_ (.A1(_04373_),
    .A2(_04403_),
    .B1(net1553),
    .Y(_00817_));
 sky130_fd_sc_hd__a211o_1 _19849_ (.A1(_02980_),
    .A2(_04347_),
    .B1(_04378_),
    .C1(_04370_),
    .X(_04405_));
 sky130_fd_sc_hd__nand2_1 _19850_ (.A(_04345_),
    .B(net928),
    .Y(_04406_));
 sky130_fd_sc_hd__o21ai_1 _19851_ (.A1(_04373_),
    .A2(_04405_),
    .B1(net929),
    .Y(_00818_));
 sky130_fd_sc_hd__and3_4 _19852_ (.A(_03207_),
    .B(_04102_),
    .C(\line_cache_idx[6] ),
    .X(_04407_));
 sky130_fd_sc_hd__nand2_1 _19853_ (.A(_04407_),
    .B(_04104_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21bo_1 _19854_ (.A1(_04408_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_8 _19855_ (.A(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _19856_ (.A0(_04101_),
    .A1(net2859),
    .S(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _19857_ (.A(_04411_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _19858_ (.A0(_04109_),
    .A1(net2528),
    .S(_04410_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _19859_ (.A(_04412_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _19860_ (.A0(_04111_),
    .A1(net2476),
    .S(_04410_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _19861_ (.A(_04413_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _19862_ (.A0(_04113_),
    .A1(net3514),
    .S(_04410_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _19863_ (.A(_04414_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _19864_ (.A0(_04115_),
    .A1(net2963),
    .S(_04410_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _19865_ (.A(_04415_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _19866_ (.A0(_04117_),
    .A1(net3488),
    .S(_04410_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _19867_ (.A(_04416_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _19868_ (.A0(_04119_),
    .A1(net3193),
    .S(_04410_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _19869_ (.A(_04417_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _19870_ (.A0(_04121_),
    .A1(net2277),
    .S(_04410_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _19871_ (.A(_04418_),
    .X(_00826_));
 sky130_fd_sc_hd__buf_4 _19872_ (.A(_04408_),
    .X(_04419_));
 sky130_fd_sc_hd__buf_4 _19873_ (.A(_03702_),
    .X(_04420_));
 sky130_fd_sc_hd__buf_4 _19874_ (.A(_04408_),
    .X(_04421_));
 sky130_fd_sc_hd__nand2_1 _19875_ (.A(_04421_),
    .B(_12185_),
    .Y(_04422_));
 sky130_fd_sc_hd__o211a_1 _19876_ (.A1(_03222_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__mux2_1 _19877_ (.A0(_04423_),
    .A1(net2985),
    .S(_04410_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _19878_ (.A(_04424_),
    .X(_00827_));
 sky130_fd_sc_hd__nand2_1 _19879_ (.A(_04421_),
    .B(_12198_),
    .Y(_04425_));
 sky130_fd_sc_hd__o211a_1 _19880_ (.A1(_03228_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_1 _19881_ (.A0(_04426_),
    .A1(net2364),
    .S(_04410_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _19882_ (.A(_04427_),
    .X(_00828_));
 sky130_fd_sc_hd__nand2_1 _19883_ (.A(_04421_),
    .B(_12206_),
    .Y(_04428_));
 sky130_fd_sc_hd__o211a_1 _19884_ (.A1(_03232_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__mux2_1 _19885_ (.A0(_04429_),
    .A1(net2609),
    .S(_04410_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _19886_ (.A(_04430_),
    .X(_00829_));
 sky130_fd_sc_hd__nand2_1 _19887_ (.A(_04421_),
    .B(_12214_),
    .Y(_04431_));
 sky130_fd_sc_hd__o211a_1 _19888_ (.A1(_03236_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__mux2_1 _19889_ (.A0(_04432_),
    .A1(net2176),
    .S(_04410_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _19890_ (.A(_04433_),
    .X(_00830_));
 sky130_fd_sc_hd__nand2_1 _19891_ (.A(_04421_),
    .B(_12222_),
    .Y(_04434_));
 sky130_fd_sc_hd__o211a_1 _19892_ (.A1(_03240_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__mux2_1 _19893_ (.A0(_04435_),
    .A1(net2637),
    .S(_04410_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _19894_ (.A(_04436_),
    .X(_00831_));
 sky130_fd_sc_hd__nand2_1 _19895_ (.A(_04421_),
    .B(_12230_),
    .Y(_04437_));
 sky130_fd_sc_hd__o211a_1 _19896_ (.A1(_03244_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__mux2_1 _19897_ (.A0(_04438_),
    .A1(net2302),
    .S(_04410_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _19898_ (.A(_04439_),
    .X(_00832_));
 sky130_fd_sc_hd__nand2_1 _19899_ (.A(_04421_),
    .B(_12238_),
    .Y(_04440_));
 sky130_fd_sc_hd__o211a_1 _19900_ (.A1(_03248_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__mux2_1 _19901_ (.A0(_04441_),
    .A1(net2428),
    .S(_04410_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _19902_ (.A(_04442_),
    .X(_00833_));
 sky130_fd_sc_hd__nand2_1 _19903_ (.A(_04421_),
    .B(_12246_),
    .Y(_04443_));
 sky130_fd_sc_hd__o211a_1 _19904_ (.A1(_03252_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__mux2_1 _19905_ (.A0(_04444_),
    .A1(net2743),
    .S(_04410_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _19906_ (.A(_04445_),
    .X(_00834_));
 sky130_fd_sc_hd__o211a_1 _19907_ (.A1(_03256_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04422_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_8 _19908_ (.A(_04409_),
    .X(_04447_));
 sky130_fd_sc_hd__mux2_1 _19909_ (.A0(_04446_),
    .A1(net2467),
    .S(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _19910_ (.A(_04448_),
    .X(_00835_));
 sky130_fd_sc_hd__o211a_1 _19911_ (.A1(_03261_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04425_),
    .X(_04449_));
 sky130_fd_sc_hd__mux2_1 _19912_ (.A0(_04449_),
    .A1(net3254),
    .S(_04447_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _19913_ (.A(_04450_),
    .X(_00836_));
 sky130_fd_sc_hd__o211a_1 _19914_ (.A1(_03264_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04428_),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(_04451_),
    .A1(net3125),
    .S(_04447_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _19916_ (.A(_04452_),
    .X(_00837_));
 sky130_fd_sc_hd__o211a_1 _19917_ (.A1(_03267_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04431_),
    .X(_04453_));
 sky130_fd_sc_hd__mux2_1 _19918_ (.A0(_04453_),
    .A1(net3112),
    .S(_04447_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _19919_ (.A(_04454_),
    .X(_00838_));
 sky130_fd_sc_hd__o211a_1 _19920_ (.A1(_03270_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04434_),
    .X(_04455_));
 sky130_fd_sc_hd__mux2_1 _19921_ (.A0(_04455_),
    .A1(net3577),
    .S(_04447_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _19922_ (.A(_04456_),
    .X(_00839_));
 sky130_fd_sc_hd__o211a_1 _19923_ (.A1(_03273_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04437_),
    .X(_04457_));
 sky130_fd_sc_hd__mux2_1 _19924_ (.A0(_04457_),
    .A1(net3184),
    .S(_04447_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _19925_ (.A(_04458_),
    .X(_00840_));
 sky130_fd_sc_hd__o211a_1 _19926_ (.A1(_03276_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04440_),
    .X(_04459_));
 sky130_fd_sc_hd__mux2_1 _19927_ (.A0(_04459_),
    .A1(net3378),
    .S(_04447_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _19928_ (.A(_04460_),
    .X(_00841_));
 sky130_fd_sc_hd__o211a_1 _19929_ (.A1(_03279_),
    .A2(_04419_),
    .B1(_04420_),
    .C1(_04443_),
    .X(_04461_));
 sky130_fd_sc_hd__mux2_1 _19930_ (.A0(_04461_),
    .A1(net2809),
    .S(_04447_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _19931_ (.A(_04462_),
    .X(_00842_));
 sky130_fd_sc_hd__buf_4 _19932_ (.A(_03702_),
    .X(_04463_));
 sky130_fd_sc_hd__o211a_1 _19933_ (.A1(_12170_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04422_),
    .X(_04464_));
 sky130_fd_sc_hd__mux2_1 _19934_ (.A0(_04464_),
    .A1(net3467),
    .S(_04447_),
    .X(_04465_));
 sky130_fd_sc_hd__clkbuf_1 _19935_ (.A(_04465_),
    .X(_00843_));
 sky130_fd_sc_hd__o211a_1 _19936_ (.A1(_12195_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04425_),
    .X(_04466_));
 sky130_fd_sc_hd__mux2_1 _19937_ (.A0(_04466_),
    .A1(net3065),
    .S(_04447_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _19938_ (.A(_04467_),
    .X(_00844_));
 sky130_fd_sc_hd__o211a_1 _19939_ (.A1(_12203_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04428_),
    .X(_04468_));
 sky130_fd_sc_hd__mux2_1 _19940_ (.A0(_04468_),
    .A1(net3491),
    .S(_04447_),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_1 _19941_ (.A(_04469_),
    .X(_00845_));
 sky130_fd_sc_hd__o211a_1 _19942_ (.A1(_12211_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04431_),
    .X(_04470_));
 sky130_fd_sc_hd__mux2_1 _19943_ (.A0(_04470_),
    .A1(net2413),
    .S(_04447_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _19944_ (.A(_04471_),
    .X(_00846_));
 sky130_fd_sc_hd__o211a_1 _19945_ (.A1(_12219_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04434_),
    .X(_04472_));
 sky130_fd_sc_hd__mux2_1 _19946_ (.A0(_04472_),
    .A1(net3622),
    .S(_04447_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _19947_ (.A(_04473_),
    .X(_00847_));
 sky130_fd_sc_hd__o211a_1 _19948_ (.A1(_12227_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04437_),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_1 _19949_ (.A0(_04474_),
    .A1(net3675),
    .S(_04447_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _19950_ (.A(_04475_),
    .X(_00848_));
 sky130_fd_sc_hd__o211a_1 _19951_ (.A1(_12235_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04440_),
    .X(_04476_));
 sky130_fd_sc_hd__mux2_1 _19952_ (.A0(_04476_),
    .A1(net3376),
    .S(_04447_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _19953_ (.A(_04477_),
    .X(_00849_));
 sky130_fd_sc_hd__o211a_1 _19954_ (.A1(_12243_),
    .A2(_04421_),
    .B1(_04463_),
    .C1(_04443_),
    .X(_04478_));
 sky130_fd_sc_hd__mux2_1 _19955_ (.A0(_04478_),
    .A1(net3569),
    .S(_04447_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _19956_ (.A(_04479_),
    .X(_00850_));
 sky130_fd_sc_hd__nand2_1 _19957_ (.A(_04407_),
    .B(_04183_),
    .Y(_04480_));
 sky130_fd_sc_hd__inv_2 _19958_ (.A(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__o21ai_4 _19959_ (.A1(_04332_),
    .A2(_04481_),
    .B1(_02818_),
    .Y(_04482_));
 sky130_fd_sc_hd__mux2_1 _19960_ (.A0(_04101_),
    .A1(net3113),
    .S(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _19961_ (.A(_04483_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _19962_ (.A0(_04109_),
    .A1(net3344),
    .S(_04482_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _19963_ (.A(_04484_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _19964_ (.A0(_04111_),
    .A1(net3219),
    .S(_04482_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _19965_ (.A(_04485_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _19966_ (.A0(_04113_),
    .A1(net2368),
    .S(_04482_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _19967_ (.A(_04486_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _19968_ (.A0(_04115_),
    .A1(net2988),
    .S(_04482_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _19969_ (.A(_04487_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _19970_ (.A0(_04117_),
    .A1(net3404),
    .S(_04482_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _19971_ (.A(_04488_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _19972_ (.A0(_04119_),
    .A1(net2960),
    .S(_04482_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _19973_ (.A(_04489_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _19974_ (.A0(_04121_),
    .A1(net3370),
    .S(_04482_),
    .X(_04490_));
 sky130_fd_sc_hd__clkbuf_1 _19975_ (.A(_04490_),
    .X(_00858_));
 sky130_fd_sc_hd__buf_4 _19976_ (.A(_04482_),
    .X(_04491_));
 sky130_fd_sc_hd__buf_4 _19977_ (.A(_04481_),
    .X(_04492_));
 sky130_fd_sc_hd__buf_4 _19978_ (.A(_04481_),
    .X(_04493_));
 sky130_fd_sc_hd__nor2_1 _19979_ (.A(_02854_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__a211o_1 _19980_ (.A1(_02852_),
    .A2(_04492_),
    .B1(_04378_),
    .C1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__buf_4 _19981_ (.A(_04482_),
    .X(_04496_));
 sky130_fd_sc_hd__nand2_1 _19982_ (.A(_04496_),
    .B(net1865),
    .Y(_04497_));
 sky130_fd_sc_hd__o21ai_1 _19983_ (.A1(_04491_),
    .A2(_04495_),
    .B1(net1866),
    .Y(_00859_));
 sky130_fd_sc_hd__nor2_1 _19984_ (.A(_02863_),
    .B(_04493_),
    .Y(_04498_));
 sky130_fd_sc_hd__a211o_1 _19985_ (.A1(_02862_),
    .A2(_04492_),
    .B1(_04378_),
    .C1(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__nand2_1 _19986_ (.A(_04496_),
    .B(net1222),
    .Y(_04500_));
 sky130_fd_sc_hd__o21ai_1 _19987_ (.A1(_04491_),
    .A2(_04499_),
    .B1(net1223),
    .Y(_00860_));
 sky130_fd_sc_hd__buf_4 _19988_ (.A(_09129_),
    .X(_04501_));
 sky130_fd_sc_hd__nor2_1 _19989_ (.A(_02870_),
    .B(_04493_),
    .Y(_04502_));
 sky130_fd_sc_hd__a211o_1 _19990_ (.A1(_02869_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__nand2_1 _19991_ (.A(_04496_),
    .B(net630),
    .Y(_04504_));
 sky130_fd_sc_hd__o21ai_1 _19992_ (.A1(_04491_),
    .A2(_04503_),
    .B1(net631),
    .Y(_00861_));
 sky130_fd_sc_hd__nor2_1 _19993_ (.A(_02877_),
    .B(_04493_),
    .Y(_04505_));
 sky130_fd_sc_hd__a211o_1 _19994_ (.A1(_02876_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__nand2_1 _19995_ (.A(_04496_),
    .B(net894),
    .Y(_04507_));
 sky130_fd_sc_hd__o21ai_1 _19996_ (.A1(_04491_),
    .A2(_04506_),
    .B1(net895),
    .Y(_00862_));
 sky130_fd_sc_hd__nor2_1 _19997_ (.A(_02884_),
    .B(_04493_),
    .Y(_04508_));
 sky130_fd_sc_hd__a211o_1 _19998_ (.A1(_02883_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__nand2_1 _19999_ (.A(_04496_),
    .B(net1008),
    .Y(_04510_));
 sky130_fd_sc_hd__o21ai_1 _20000_ (.A1(_04491_),
    .A2(_04509_),
    .B1(net1009),
    .Y(_00863_));
 sky130_fd_sc_hd__nor2_1 _20001_ (.A(_02891_),
    .B(_04493_),
    .Y(_04511_));
 sky130_fd_sc_hd__a211o_1 _20002_ (.A1(_02890_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__nand2_1 _20003_ (.A(_04496_),
    .B(net1606),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ai_1 _20004_ (.A1(_04491_),
    .A2(_04512_),
    .B1(net1607),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_1 _20005_ (.A(_02898_),
    .B(_04493_),
    .Y(_04514_));
 sky130_fd_sc_hd__a211o_1 _20006_ (.A1(_02897_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__nand2_1 _20007_ (.A(_04496_),
    .B(net1556),
    .Y(_04516_));
 sky130_fd_sc_hd__o21ai_1 _20008_ (.A1(_04491_),
    .A2(_04515_),
    .B1(net1557),
    .Y(_00865_));
 sky130_fd_sc_hd__nor2_1 _20009_ (.A(_02905_),
    .B(_04493_),
    .Y(_04517_));
 sky130_fd_sc_hd__a211o_1 _20010_ (.A1(_02904_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _20011_ (.A(_04496_),
    .B(net992),
    .Y(_04519_));
 sky130_fd_sc_hd__o21ai_1 _20012_ (.A1(_04491_),
    .A2(_04518_),
    .B1(net993),
    .Y(_00866_));
 sky130_fd_sc_hd__buf_4 _20013_ (.A(_04482_),
    .X(_04520_));
 sky130_fd_sc_hd__a211o_1 _20014_ (.A1(_02912_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04494_),
    .X(_04521_));
 sky130_fd_sc_hd__nand2_1 _20015_ (.A(_04496_),
    .B(net1875),
    .Y(_04522_));
 sky130_fd_sc_hd__o21ai_1 _20016_ (.A1(_04520_),
    .A2(_04521_),
    .B1(net1876),
    .Y(_00867_));
 sky130_fd_sc_hd__a211o_1 _20017_ (.A1(_02917_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04498_),
    .X(_04523_));
 sky130_fd_sc_hd__nand2_1 _20018_ (.A(_04496_),
    .B(net614),
    .Y(_04524_));
 sky130_fd_sc_hd__o21ai_1 _20019_ (.A1(_04520_),
    .A2(_04523_),
    .B1(net615),
    .Y(_00868_));
 sky130_fd_sc_hd__a211o_1 _20020_ (.A1(_02922_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04502_),
    .X(_04525_));
 sky130_fd_sc_hd__nand2_1 _20021_ (.A(_04496_),
    .B(net612),
    .Y(_04526_));
 sky130_fd_sc_hd__o21ai_1 _20022_ (.A1(_04520_),
    .A2(_04525_),
    .B1(net613),
    .Y(_00869_));
 sky130_fd_sc_hd__a211o_1 _20023_ (.A1(_02928_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04505_),
    .X(_04527_));
 sky130_fd_sc_hd__nand2_1 _20024_ (.A(_04496_),
    .B(net1310),
    .Y(_04528_));
 sky130_fd_sc_hd__o21ai_1 _20025_ (.A1(_04520_),
    .A2(_04527_),
    .B1(net1311),
    .Y(_00870_));
 sky130_fd_sc_hd__a211o_1 _20026_ (.A1(_02933_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04508_),
    .X(_04529_));
 sky130_fd_sc_hd__nand2_1 _20027_ (.A(_04496_),
    .B(net972),
    .Y(_04530_));
 sky130_fd_sc_hd__o21ai_1 _20028_ (.A1(_04520_),
    .A2(_04529_),
    .B1(net973),
    .Y(_00871_));
 sky130_fd_sc_hd__a211o_1 _20029_ (.A1(_02938_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04511_),
    .X(_04531_));
 sky130_fd_sc_hd__nand2_1 _20030_ (.A(_04496_),
    .B(net1526),
    .Y(_04532_));
 sky130_fd_sc_hd__o21ai_1 _20031_ (.A1(_04520_),
    .A2(_04531_),
    .B1(net1527),
    .Y(_00872_));
 sky130_fd_sc_hd__a211o_1 _20032_ (.A1(_02943_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04514_),
    .X(_04533_));
 sky130_fd_sc_hd__nand2_1 _20033_ (.A(_04496_),
    .B(net1522),
    .Y(_04534_));
 sky130_fd_sc_hd__o21ai_1 _20034_ (.A1(_04520_),
    .A2(_04533_),
    .B1(net1523),
    .Y(_00873_));
 sky130_fd_sc_hd__a211o_1 _20035_ (.A1(_02948_),
    .A2(_04492_),
    .B1(_04501_),
    .C1(_04517_),
    .X(_04535_));
 sky130_fd_sc_hd__nand2_1 _20036_ (.A(_04496_),
    .B(net1378),
    .Y(_04536_));
 sky130_fd_sc_hd__o21ai_1 _20037_ (.A1(_04520_),
    .A2(_04535_),
    .B1(net1379),
    .Y(_00874_));
 sky130_fd_sc_hd__a211o_1 _20038_ (.A1(_02952_),
    .A2(_04493_),
    .B1(_04501_),
    .C1(_04494_),
    .X(_04537_));
 sky130_fd_sc_hd__nand2_1 _20039_ (.A(_04491_),
    .B(net1102),
    .Y(_04538_));
 sky130_fd_sc_hd__o21ai_1 _20040_ (.A1(_04520_),
    .A2(_04537_),
    .B1(net1103),
    .Y(_00875_));
 sky130_fd_sc_hd__a211o_1 _20041_ (.A1(_02956_),
    .A2(_04493_),
    .B1(_04501_),
    .C1(_04498_),
    .X(_04539_));
 sky130_fd_sc_hd__nand2_1 _20042_ (.A(_04491_),
    .B(net1442),
    .Y(_04540_));
 sky130_fd_sc_hd__o21ai_1 _20043_ (.A1(_04520_),
    .A2(_04539_),
    .B1(net1443),
    .Y(_00876_));
 sky130_fd_sc_hd__clkbuf_8 _20044_ (.A(_09129_),
    .X(_04541_));
 sky130_fd_sc_hd__a211o_1 _20045_ (.A1(_02960_),
    .A2(_04493_),
    .B1(_04541_),
    .C1(_04502_),
    .X(_04542_));
 sky130_fd_sc_hd__nand2_1 _20046_ (.A(_04491_),
    .B(net1042),
    .Y(_04543_));
 sky130_fd_sc_hd__o21ai_1 _20047_ (.A1(_04520_),
    .A2(_04542_),
    .B1(net1043),
    .Y(_00877_));
 sky130_fd_sc_hd__a211o_1 _20048_ (.A1(_02964_),
    .A2(_04493_),
    .B1(_04541_),
    .C1(_04505_),
    .X(_04544_));
 sky130_fd_sc_hd__nand2_1 _20049_ (.A(_04491_),
    .B(net848),
    .Y(_04545_));
 sky130_fd_sc_hd__o21ai_1 _20050_ (.A1(_04520_),
    .A2(_04544_),
    .B1(net849),
    .Y(_00878_));
 sky130_fd_sc_hd__a211o_1 _20051_ (.A1(_02968_),
    .A2(_04493_),
    .B1(_04541_),
    .C1(_04508_),
    .X(_04546_));
 sky130_fd_sc_hd__nand2_1 _20052_ (.A(_04491_),
    .B(net884),
    .Y(_04547_));
 sky130_fd_sc_hd__o21ai_1 _20053_ (.A1(_04520_),
    .A2(_04546_),
    .B1(net885),
    .Y(_00879_));
 sky130_fd_sc_hd__a211o_1 _20054_ (.A1(_02972_),
    .A2(_04493_),
    .B1(_04541_),
    .C1(_04511_),
    .X(_04548_));
 sky130_fd_sc_hd__nand2_1 _20055_ (.A(_04491_),
    .B(net662),
    .Y(_04549_));
 sky130_fd_sc_hd__o21ai_1 _20056_ (.A1(_04520_),
    .A2(_04548_),
    .B1(net663),
    .Y(_00880_));
 sky130_fd_sc_hd__a211o_1 _20057_ (.A1(_02976_),
    .A2(_04493_),
    .B1(_04541_),
    .C1(_04514_),
    .X(_04550_));
 sky130_fd_sc_hd__nand2_1 _20058_ (.A(_04491_),
    .B(net874),
    .Y(_04551_));
 sky130_fd_sc_hd__o21ai_1 _20059_ (.A1(_04520_),
    .A2(_04550_),
    .B1(net875),
    .Y(_00881_));
 sky130_fd_sc_hd__a211o_1 _20060_ (.A1(_02980_),
    .A2(_04493_),
    .B1(_04541_),
    .C1(_04517_),
    .X(_04552_));
 sky130_fd_sc_hd__nand2_1 _20061_ (.A(_04491_),
    .B(net1216),
    .Y(_04553_));
 sky130_fd_sc_hd__o21ai_1 _20062_ (.A1(_04520_),
    .A2(_04552_),
    .B1(net1217),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _20063_ (.A(_04407_),
    .B(_04257_),
    .Y(_04554_));
 sky130_fd_sc_hd__inv_2 _20064_ (.A(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__o21ai_4 _20065_ (.A1(_04332_),
    .A2(_04555_),
    .B1(_02818_),
    .Y(_04556_));
 sky130_fd_sc_hd__mux2_1 _20066_ (.A0(_04101_),
    .A1(net2900),
    .S(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_1 _20067_ (.A(_04557_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _20068_ (.A0(_04109_),
    .A1(net2702),
    .S(_04556_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _20069_ (.A(_04558_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _20070_ (.A0(_04111_),
    .A1(net2148),
    .S(_04556_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _20071_ (.A(_04559_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _20072_ (.A0(_04113_),
    .A1(net3526),
    .S(_04556_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _20073_ (.A(_04560_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _20074_ (.A0(_04115_),
    .A1(net2234),
    .S(_04556_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _20075_ (.A(_04561_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _20076_ (.A0(_04117_),
    .A1(net3267),
    .S(_04556_),
    .X(_04562_));
 sky130_fd_sc_hd__clkbuf_1 _20077_ (.A(_04562_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _20078_ (.A0(_04119_),
    .A1(net2384),
    .S(_04556_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _20079_ (.A(_04563_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _20080_ (.A0(_04121_),
    .A1(net3036),
    .S(_04556_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _20081_ (.A(_04564_),
    .X(_00890_));
 sky130_fd_sc_hd__buf_4 _20082_ (.A(_04556_),
    .X(_04565_));
 sky130_fd_sc_hd__buf_4 _20083_ (.A(_04555_),
    .X(_04566_));
 sky130_fd_sc_hd__buf_4 _20084_ (.A(_04555_),
    .X(_04567_));
 sky130_fd_sc_hd__nor2_1 _20085_ (.A(_02854_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__a211o_1 _20086_ (.A1(_02852_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__buf_4 _20087_ (.A(_04556_),
    .X(_04570_));
 sky130_fd_sc_hd__nand2_1 _20088_ (.A(_04570_),
    .B(net864),
    .Y(_04571_));
 sky130_fd_sc_hd__o21ai_1 _20089_ (.A1(_04565_),
    .A2(_04569_),
    .B1(net865),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2_1 _20090_ (.A(_02863_),
    .B(_04567_),
    .Y(_04572_));
 sky130_fd_sc_hd__a211o_1 _20091_ (.A1(_02862_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__nand2_1 _20092_ (.A(_04570_),
    .B(net734),
    .Y(_04574_));
 sky130_fd_sc_hd__o21ai_1 _20093_ (.A1(_04565_),
    .A2(_04573_),
    .B1(net735),
    .Y(_00892_));
 sky130_fd_sc_hd__nor2_1 _20094_ (.A(_02870_),
    .B(_04567_),
    .Y(_04575_));
 sky130_fd_sc_hd__a211o_1 _20095_ (.A1(_02869_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__nand2_1 _20096_ (.A(_04570_),
    .B(net620),
    .Y(_04577_));
 sky130_fd_sc_hd__o21ai_1 _20097_ (.A1(_04565_),
    .A2(_04576_),
    .B1(net621),
    .Y(_00893_));
 sky130_fd_sc_hd__nor2_1 _20098_ (.A(_02877_),
    .B(_04567_),
    .Y(_04578_));
 sky130_fd_sc_hd__a211o_1 _20099_ (.A1(_02876_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__nand2_1 _20100_ (.A(_04570_),
    .B(net700),
    .Y(_04580_));
 sky130_fd_sc_hd__o21ai_1 _20101_ (.A1(_04565_),
    .A2(_04579_),
    .B1(net701),
    .Y(_00894_));
 sky130_fd_sc_hd__nor2_1 _20102_ (.A(_02884_),
    .B(_04567_),
    .Y(_04581_));
 sky130_fd_sc_hd__a211o_1 _20103_ (.A1(_02883_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _20104_ (.A(_04570_),
    .B(net1618),
    .Y(_04583_));
 sky130_fd_sc_hd__o21ai_1 _20105_ (.A1(_04565_),
    .A2(_04582_),
    .B1(net1619),
    .Y(_00895_));
 sky130_fd_sc_hd__nor2_1 _20106_ (.A(_02891_),
    .B(_04567_),
    .Y(_04584_));
 sky130_fd_sc_hd__a211o_1 _20107_ (.A1(_02890_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__nand2_1 _20108_ (.A(_04570_),
    .B(net1448),
    .Y(_04586_));
 sky130_fd_sc_hd__o21ai_1 _20109_ (.A1(_04565_),
    .A2(_04585_),
    .B1(net1449),
    .Y(_00896_));
 sky130_fd_sc_hd__nor2_1 _20110_ (.A(_02898_),
    .B(_04567_),
    .Y(_04587_));
 sky130_fd_sc_hd__a211o_1 _20111_ (.A1(_02897_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__nand2_1 _20112_ (.A(_04570_),
    .B(net774),
    .Y(_04589_));
 sky130_fd_sc_hd__o21ai_1 _20113_ (.A1(_04565_),
    .A2(_04588_),
    .B1(net775),
    .Y(_00897_));
 sky130_fd_sc_hd__nor2_1 _20114_ (.A(_02905_),
    .B(_04567_),
    .Y(_04590_));
 sky130_fd_sc_hd__a211o_1 _20115_ (.A1(_02904_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_1 _20116_ (.A(_04570_),
    .B(net1156),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_1 _20117_ (.A1(_04565_),
    .A2(_04591_),
    .B1(net1157),
    .Y(_00898_));
 sky130_fd_sc_hd__buf_4 _20118_ (.A(_04556_),
    .X(_04593_));
 sky130_fd_sc_hd__a211o_1 _20119_ (.A1(_02912_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04568_),
    .X(_04594_));
 sky130_fd_sc_hd__nand2_1 _20120_ (.A(_04570_),
    .B(net1939),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_1 _20121_ (.A1(_04593_),
    .A2(_04594_),
    .B1(_04595_),
    .Y(_00899_));
 sky130_fd_sc_hd__a211o_1 _20122_ (.A1(_02917_),
    .A2(_04566_),
    .B1(_04541_),
    .C1(_04572_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_1 _20123_ (.A(_04570_),
    .B(net1436),
    .Y(_04597_));
 sky130_fd_sc_hd__o21ai_1 _20124_ (.A1(_04593_),
    .A2(_04596_),
    .B1(net1437),
    .Y(_00900_));
 sky130_fd_sc_hd__buf_8 _20125_ (.A(_09057_),
    .X(_04598_));
 sky130_fd_sc_hd__buf_4 _20126_ (.A(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__a211o_1 _20127_ (.A1(_02922_),
    .A2(_04566_),
    .B1(_04599_),
    .C1(_04575_),
    .X(_04600_));
 sky130_fd_sc_hd__nand2_1 _20128_ (.A(_04570_),
    .B(net1344),
    .Y(_04601_));
 sky130_fd_sc_hd__o21ai_1 _20129_ (.A1(_04593_),
    .A2(_04600_),
    .B1(net1345),
    .Y(_00901_));
 sky130_fd_sc_hd__a211o_1 _20130_ (.A1(_02928_),
    .A2(_04566_),
    .B1(_04599_),
    .C1(_04578_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_1 _20131_ (.A(_04570_),
    .B(net1278),
    .Y(_04603_));
 sky130_fd_sc_hd__o21ai_1 _20132_ (.A1(_04593_),
    .A2(_04602_),
    .B1(net1279),
    .Y(_00902_));
 sky130_fd_sc_hd__a211o_1 _20133_ (.A1(_02933_),
    .A2(_04566_),
    .B1(_04599_),
    .C1(_04581_),
    .X(_04604_));
 sky130_fd_sc_hd__nand2_1 _20134_ (.A(_04570_),
    .B(net1662),
    .Y(_04605_));
 sky130_fd_sc_hd__o21ai_1 _20135_ (.A1(_04593_),
    .A2(_04604_),
    .B1(net1663),
    .Y(_00903_));
 sky130_fd_sc_hd__a211o_1 _20136_ (.A1(_02938_),
    .A2(_04566_),
    .B1(_04599_),
    .C1(_04584_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2_1 _20137_ (.A(_04570_),
    .B(net766),
    .Y(_04607_));
 sky130_fd_sc_hd__o21ai_1 _20138_ (.A1(_04593_),
    .A2(_04606_),
    .B1(net767),
    .Y(_00904_));
 sky130_fd_sc_hd__a211o_1 _20139_ (.A1(_02943_),
    .A2(_04566_),
    .B1(_04599_),
    .C1(_04587_),
    .X(_04608_));
 sky130_fd_sc_hd__nand2_1 _20140_ (.A(_04570_),
    .B(net1426),
    .Y(_04609_));
 sky130_fd_sc_hd__o21ai_1 _20141_ (.A1(_04593_),
    .A2(_04608_),
    .B1(net1427),
    .Y(_00905_));
 sky130_fd_sc_hd__a211o_1 _20142_ (.A1(_02948_),
    .A2(_04566_),
    .B1(_04599_),
    .C1(_04590_),
    .X(_04610_));
 sky130_fd_sc_hd__nand2_1 _20143_ (.A(_04570_),
    .B(net698),
    .Y(_04611_));
 sky130_fd_sc_hd__o21ai_1 _20144_ (.A1(_04593_),
    .A2(_04610_),
    .B1(net699),
    .Y(_00906_));
 sky130_fd_sc_hd__a211o_1 _20145_ (.A1(_02952_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04568_),
    .X(_04612_));
 sky130_fd_sc_hd__nand2_1 _20146_ (.A(_04565_),
    .B(net1414),
    .Y(_04613_));
 sky130_fd_sc_hd__o21ai_1 _20147_ (.A1(_04593_),
    .A2(_04612_),
    .B1(net1415),
    .Y(_00907_));
 sky130_fd_sc_hd__a211o_1 _20148_ (.A1(_02956_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04572_),
    .X(_04614_));
 sky130_fd_sc_hd__nand2_1 _20149_ (.A(_04565_),
    .B(net1160),
    .Y(_04615_));
 sky130_fd_sc_hd__o21ai_1 _20150_ (.A1(_04593_),
    .A2(_04614_),
    .B1(net1161),
    .Y(_00908_));
 sky130_fd_sc_hd__a211o_1 _20151_ (.A1(_02960_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04575_),
    .X(_04616_));
 sky130_fd_sc_hd__nand2_1 _20152_ (.A(_04565_),
    .B(net820),
    .Y(_04617_));
 sky130_fd_sc_hd__o21ai_1 _20153_ (.A1(_04593_),
    .A2(_04616_),
    .B1(net821),
    .Y(_00909_));
 sky130_fd_sc_hd__a211o_1 _20154_ (.A1(_02964_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04578_),
    .X(_04618_));
 sky130_fd_sc_hd__nand2_1 _20155_ (.A(_04565_),
    .B(net748),
    .Y(_04619_));
 sky130_fd_sc_hd__o21ai_1 _20156_ (.A1(_04593_),
    .A2(_04618_),
    .B1(net749),
    .Y(_00910_));
 sky130_fd_sc_hd__a211o_1 _20157_ (.A1(_02968_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04581_),
    .X(_04620_));
 sky130_fd_sc_hd__nand2_1 _20158_ (.A(_04565_),
    .B(net1014),
    .Y(_04621_));
 sky130_fd_sc_hd__o21ai_1 _20159_ (.A1(_04593_),
    .A2(_04620_),
    .B1(net1015),
    .Y(_00911_));
 sky130_fd_sc_hd__a211o_1 _20160_ (.A1(_02972_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04584_),
    .X(_04622_));
 sky130_fd_sc_hd__nand2_1 _20161_ (.A(_04565_),
    .B(net672),
    .Y(_04623_));
 sky130_fd_sc_hd__o21ai_1 _20162_ (.A1(_04593_),
    .A2(_04622_),
    .B1(net673),
    .Y(_00912_));
 sky130_fd_sc_hd__a211o_1 _20163_ (.A1(_02976_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04587_),
    .X(_04624_));
 sky130_fd_sc_hd__nand2_1 _20164_ (.A(_04565_),
    .B(net1400),
    .Y(_04625_));
 sky130_fd_sc_hd__o21ai_1 _20165_ (.A1(_04593_),
    .A2(_04624_),
    .B1(net1401),
    .Y(_00913_));
 sky130_fd_sc_hd__a211o_1 _20166_ (.A1(_02980_),
    .A2(_04567_),
    .B1(_04599_),
    .C1(_04590_),
    .X(_04626_));
 sky130_fd_sc_hd__nand2_1 _20167_ (.A(_04565_),
    .B(net1570),
    .Y(_04627_));
 sky130_fd_sc_hd__o21ai_1 _20168_ (.A1(_04593_),
    .A2(_04626_),
    .B1(net1571),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _20169_ (.A(_04407_),
    .B(_04333_),
    .Y(_04628_));
 sky130_fd_sc_hd__inv_2 _20170_ (.A(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__o21ai_4 _20171_ (.A1(_04332_),
    .A2(_04629_),
    .B1(_02818_),
    .Y(_04630_));
 sky130_fd_sc_hd__mux2_1 _20172_ (.A0(_04101_),
    .A1(net2316),
    .S(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_1 _20173_ (.A(_04631_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _20174_ (.A0(_04109_),
    .A1(net2808),
    .S(_04630_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _20175_ (.A(_04632_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _20176_ (.A0(_04111_),
    .A1(net3532),
    .S(_04630_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _20177_ (.A(_04633_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _20178_ (.A0(_04113_),
    .A1(net3730),
    .S(_04630_),
    .X(_04634_));
 sky130_fd_sc_hd__clkbuf_1 _20179_ (.A(_04634_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _20180_ (.A0(_04115_),
    .A1(net3026),
    .S(_04630_),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _20181_ (.A(_04635_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _20182_ (.A0(_04117_),
    .A1(net3654),
    .S(_04630_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _20183_ (.A(_04636_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _20184_ (.A0(_04119_),
    .A1(net2228),
    .S(_04630_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_1 _20185_ (.A(_04637_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _20186_ (.A0(_04121_),
    .A1(net2186),
    .S(_04630_),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _20187_ (.A(_04638_),
    .X(_00922_));
 sky130_fd_sc_hd__buf_4 _20188_ (.A(_04630_),
    .X(_04639_));
 sky130_fd_sc_hd__buf_4 _20189_ (.A(_04629_),
    .X(_04640_));
 sky130_fd_sc_hd__buf_4 _20190_ (.A(_04629_),
    .X(_04641_));
 sky130_fd_sc_hd__nor2_1 _20191_ (.A(_02854_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__a211o_1 _20192_ (.A1(_02852_),
    .A2(_04640_),
    .B1(_04599_),
    .C1(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__buf_4 _20193_ (.A(_04630_),
    .X(_04644_));
 sky130_fd_sc_hd__nand2_1 _20194_ (.A(_04644_),
    .B(net770),
    .Y(_04645_));
 sky130_fd_sc_hd__o21ai_1 _20195_ (.A1(_04639_),
    .A2(_04643_),
    .B1(net771),
    .Y(_00923_));
 sky130_fd_sc_hd__nor2_1 _20196_ (.A(_02863_),
    .B(_04641_),
    .Y(_04646_));
 sky130_fd_sc_hd__a211o_1 _20197_ (.A1(_02862_),
    .A2(_04640_),
    .B1(_04599_),
    .C1(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__nand2_1 _20198_ (.A(_04644_),
    .B(net544),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ai_1 _20199_ (.A1(_04639_),
    .A2(_04647_),
    .B1(net545),
    .Y(_00924_));
 sky130_fd_sc_hd__buf_4 _20200_ (.A(_04598_),
    .X(_04649_));
 sky130_fd_sc_hd__nor2_1 _20201_ (.A(_02870_),
    .B(_04641_),
    .Y(_04650_));
 sky130_fd_sc_hd__a211o_1 _20202_ (.A1(_02869_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__nand2_1 _20203_ (.A(_04644_),
    .B(net642),
    .Y(_04652_));
 sky130_fd_sc_hd__o21ai_1 _20204_ (.A1(_04639_),
    .A2(_04651_),
    .B1(net643),
    .Y(_00925_));
 sky130_fd_sc_hd__nor2_1 _20205_ (.A(_02877_),
    .B(_04641_),
    .Y(_04653_));
 sky130_fd_sc_hd__a211o_1 _20206_ (.A1(_02876_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__nand2_1 _20207_ (.A(_04644_),
    .B(net718),
    .Y(_04655_));
 sky130_fd_sc_hd__o21ai_1 _20208_ (.A1(_04639_),
    .A2(_04654_),
    .B1(net719),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_1 _20209_ (.A(_02884_),
    .B(_04641_),
    .Y(_04656_));
 sky130_fd_sc_hd__a211o_1 _20210_ (.A1(_02883_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _20211_ (.A(_04644_),
    .B(net654),
    .Y(_04658_));
 sky130_fd_sc_hd__o21ai_1 _20212_ (.A1(_04639_),
    .A2(_04657_),
    .B1(net655),
    .Y(_00927_));
 sky130_fd_sc_hd__nor2_1 _20213_ (.A(_02891_),
    .B(_04641_),
    .Y(_04659_));
 sky130_fd_sc_hd__a211o_1 _20214_ (.A1(_02890_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__nand2_1 _20215_ (.A(_04644_),
    .B(net776),
    .Y(_04661_));
 sky130_fd_sc_hd__o21ai_1 _20216_ (.A1(_04639_),
    .A2(_04660_),
    .B1(net777),
    .Y(_00928_));
 sky130_fd_sc_hd__nor2_1 _20217_ (.A(_02898_),
    .B(_04641_),
    .Y(_04662_));
 sky130_fd_sc_hd__a211o_1 _20218_ (.A1(_02897_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__nand2_1 _20219_ (.A(_04644_),
    .B(net1590),
    .Y(_04664_));
 sky130_fd_sc_hd__o21ai_1 _20220_ (.A1(_04639_),
    .A2(_04663_),
    .B1(net1591),
    .Y(_00929_));
 sky130_fd_sc_hd__nor2_1 _20221_ (.A(_02905_),
    .B(_04641_),
    .Y(_04665_));
 sky130_fd_sc_hd__a211o_1 _20222_ (.A1(_02904_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__nand2_1 _20223_ (.A(_04644_),
    .B(net978),
    .Y(_04667_));
 sky130_fd_sc_hd__o21ai_1 _20224_ (.A1(_04639_),
    .A2(_04666_),
    .B1(net979),
    .Y(_00930_));
 sky130_fd_sc_hd__buf_4 _20225_ (.A(_04630_),
    .X(_04668_));
 sky130_fd_sc_hd__a211o_1 _20226_ (.A1(_02912_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04642_),
    .X(_04669_));
 sky130_fd_sc_hd__nand2_1 _20227_ (.A(_04644_),
    .B(net1474),
    .Y(_04670_));
 sky130_fd_sc_hd__o21ai_1 _20228_ (.A1(_04668_),
    .A2(_04669_),
    .B1(net1475),
    .Y(_00931_));
 sky130_fd_sc_hd__a211o_1 _20229_ (.A1(_02917_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04646_),
    .X(_04671_));
 sky130_fd_sc_hd__nand2_1 _20230_ (.A(_04644_),
    .B(net882),
    .Y(_04672_));
 sky130_fd_sc_hd__o21ai_1 _20231_ (.A1(_04668_),
    .A2(_04671_),
    .B1(net883),
    .Y(_00932_));
 sky130_fd_sc_hd__a211o_1 _20232_ (.A1(_02922_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04650_),
    .X(_04673_));
 sky130_fd_sc_hd__nand2_1 _20233_ (.A(_04644_),
    .B(net720),
    .Y(_04674_));
 sky130_fd_sc_hd__o21ai_1 _20234_ (.A1(_04668_),
    .A2(_04673_),
    .B1(net721),
    .Y(_00933_));
 sky130_fd_sc_hd__a211o_1 _20235_ (.A1(_02928_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04653_),
    .X(_04675_));
 sky130_fd_sc_hd__nand2_1 _20236_ (.A(_04644_),
    .B(net1054),
    .Y(_04676_));
 sky130_fd_sc_hd__o21ai_1 _20237_ (.A1(_04668_),
    .A2(_04675_),
    .B1(net1055),
    .Y(_00934_));
 sky130_fd_sc_hd__a211o_1 _20238_ (.A1(_02933_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04656_),
    .X(_04677_));
 sky130_fd_sc_hd__nand2_1 _20239_ (.A(_04644_),
    .B(net1374),
    .Y(_04678_));
 sky130_fd_sc_hd__o21ai_1 _20240_ (.A1(_04668_),
    .A2(_04677_),
    .B1(net1375),
    .Y(_00935_));
 sky130_fd_sc_hd__a211o_1 _20241_ (.A1(_02938_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04659_),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _20242_ (.A(_04644_),
    .B(net1889),
    .Y(_04680_));
 sky130_fd_sc_hd__o21ai_1 _20243_ (.A1(_04668_),
    .A2(_04679_),
    .B1(net1890),
    .Y(_00936_));
 sky130_fd_sc_hd__a211o_1 _20244_ (.A1(_02943_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04662_),
    .X(_04681_));
 sky130_fd_sc_hd__nand2_1 _20245_ (.A(_04644_),
    .B(net1416),
    .Y(_04682_));
 sky130_fd_sc_hd__o21ai_1 _20246_ (.A1(_04668_),
    .A2(_04681_),
    .B1(net1417),
    .Y(_00937_));
 sky130_fd_sc_hd__a211o_1 _20247_ (.A1(_02948_),
    .A2(_04640_),
    .B1(_04649_),
    .C1(_04665_),
    .X(_04683_));
 sky130_fd_sc_hd__nand2_1 _20248_ (.A(_04644_),
    .B(net1300),
    .Y(_04684_));
 sky130_fd_sc_hd__o21ai_1 _20249_ (.A1(_04668_),
    .A2(_04683_),
    .B1(net1301),
    .Y(_00938_));
 sky130_fd_sc_hd__a211o_1 _20250_ (.A1(_02952_),
    .A2(_04641_),
    .B1(_04649_),
    .C1(_04642_),
    .X(_04685_));
 sky130_fd_sc_hd__nand2_1 _20251_ (.A(_04639_),
    .B(net1566),
    .Y(_04686_));
 sky130_fd_sc_hd__o21ai_1 _20252_ (.A1(_04668_),
    .A2(_04685_),
    .B1(net1567),
    .Y(_00939_));
 sky130_fd_sc_hd__a211o_1 _20253_ (.A1(_02956_),
    .A2(_04641_),
    .B1(_04649_),
    .C1(_04646_),
    .X(_04687_));
 sky130_fd_sc_hd__nand2_1 _20254_ (.A(_04639_),
    .B(net982),
    .Y(_04688_));
 sky130_fd_sc_hd__o21ai_1 _20255_ (.A1(_04668_),
    .A2(_04687_),
    .B1(net983),
    .Y(_00940_));
 sky130_fd_sc_hd__clkbuf_8 _20256_ (.A(_04598_),
    .X(_04689_));
 sky130_fd_sc_hd__a211o_1 _20257_ (.A1(_02960_),
    .A2(_04641_),
    .B1(_04689_),
    .C1(_04650_),
    .X(_04690_));
 sky130_fd_sc_hd__nand2_1 _20258_ (.A(_04639_),
    .B(net1660),
    .Y(_04691_));
 sky130_fd_sc_hd__o21ai_1 _20259_ (.A1(_04668_),
    .A2(_04690_),
    .B1(net1661),
    .Y(_00941_));
 sky130_fd_sc_hd__a211o_1 _20260_ (.A1(_02964_),
    .A2(_04641_),
    .B1(_04689_),
    .C1(_04653_),
    .X(_04692_));
 sky130_fd_sc_hd__nand2_1 _20261_ (.A(_04639_),
    .B(net1198),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ai_1 _20262_ (.A1(_04668_),
    .A2(_04692_),
    .B1(net1199),
    .Y(_00942_));
 sky130_fd_sc_hd__a211o_1 _20263_ (.A1(_02968_),
    .A2(_04641_),
    .B1(_04689_),
    .C1(_04656_),
    .X(_04694_));
 sky130_fd_sc_hd__nand2_1 _20264_ (.A(_04639_),
    .B(net1564),
    .Y(_04695_));
 sky130_fd_sc_hd__o21ai_1 _20265_ (.A1(_04668_),
    .A2(_04694_),
    .B1(net1565),
    .Y(_00943_));
 sky130_fd_sc_hd__a211o_1 _20266_ (.A1(_02972_),
    .A2(_04641_),
    .B1(_04689_),
    .C1(_04659_),
    .X(_04696_));
 sky130_fd_sc_hd__nand2_1 _20267_ (.A(_04639_),
    .B(net790),
    .Y(_04697_));
 sky130_fd_sc_hd__o21ai_1 _20268_ (.A1(_04668_),
    .A2(_04696_),
    .B1(net791),
    .Y(_00944_));
 sky130_fd_sc_hd__a211o_1 _20269_ (.A1(_02976_),
    .A2(_04641_),
    .B1(_04689_),
    .C1(_04662_),
    .X(_04698_));
 sky130_fd_sc_hd__nand2_1 _20270_ (.A(_04639_),
    .B(net652),
    .Y(_04699_));
 sky130_fd_sc_hd__o21ai_1 _20271_ (.A1(_04668_),
    .A2(_04698_),
    .B1(net653),
    .Y(_00945_));
 sky130_fd_sc_hd__a211o_1 _20272_ (.A1(_02980_),
    .A2(_04641_),
    .B1(_04689_),
    .C1(_04665_),
    .X(_04700_));
 sky130_fd_sc_hd__nand2_1 _20273_ (.A(_04639_),
    .B(net754),
    .Y(_04701_));
 sky130_fd_sc_hd__o21ai_1 _20274_ (.A1(_04668_),
    .A2(_04700_),
    .B1(net755),
    .Y(_00946_));
 sky130_fd_sc_hd__and3_4 _20275_ (.A(_03516_),
    .B(_04102_),
    .C(\line_cache_idx[6] ),
    .X(_04702_));
 sky130_fd_sc_hd__nand2_1 _20276_ (.A(_04702_),
    .B(_04104_),
    .Y(_04703_));
 sky130_fd_sc_hd__a21bo_1 _20277_ (.A1(_04703_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_04704_));
 sky130_fd_sc_hd__buf_6 _20278_ (.A(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__mux2_1 _20279_ (.A0(_04101_),
    .A1(net3290),
    .S(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__clkbuf_1 _20280_ (.A(_04706_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _20281_ (.A0(_04109_),
    .A1(net2341),
    .S(_04705_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _20282_ (.A(_04707_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _20283_ (.A0(_04111_),
    .A1(net3610),
    .S(_04705_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_1 _20284_ (.A(_04708_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _20285_ (.A0(_04113_),
    .A1(net2650),
    .S(_04705_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _20286_ (.A(_04709_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _20287_ (.A0(_04115_),
    .A1(net2844),
    .S(_04705_),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_1 _20288_ (.A(_04710_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _20289_ (.A0(_04117_),
    .A1(net3301),
    .S(_04705_),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _20290_ (.A(_04711_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _20291_ (.A0(_04119_),
    .A1(net2181),
    .S(_04705_),
    .X(_04712_));
 sky130_fd_sc_hd__clkbuf_1 _20292_ (.A(_04712_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _20293_ (.A0(_04121_),
    .A1(net2548),
    .S(_04705_),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _20294_ (.A(_04713_),
    .X(_00954_));
 sky130_fd_sc_hd__buf_4 _20295_ (.A(_04703_),
    .X(_04714_));
 sky130_fd_sc_hd__buf_4 _20296_ (.A(_04703_),
    .X(_04715_));
 sky130_fd_sc_hd__nand2_1 _20297_ (.A(_04715_),
    .B(_12185_),
    .Y(_04716_));
 sky130_fd_sc_hd__o211a_1 _20298_ (.A1(_03222_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__mux2_1 _20299_ (.A0(_04717_),
    .A1(net2425),
    .S(_04705_),
    .X(_04718_));
 sky130_fd_sc_hd__clkbuf_1 _20300_ (.A(_04718_),
    .X(_00955_));
 sky130_fd_sc_hd__nand2_1 _20301_ (.A(_04715_),
    .B(_12198_),
    .Y(_04719_));
 sky130_fd_sc_hd__o211a_1 _20302_ (.A1(_03228_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__mux2_1 _20303_ (.A0(_04720_),
    .A1(net3264),
    .S(_04705_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_1 _20304_ (.A(_04721_),
    .X(_00956_));
 sky130_fd_sc_hd__nand2_1 _20305_ (.A(_04715_),
    .B(_12206_),
    .Y(_04722_));
 sky130_fd_sc_hd__o211a_1 _20306_ (.A1(_03232_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__mux2_1 _20307_ (.A0(_04723_),
    .A1(net3153),
    .S(_04705_),
    .X(_04724_));
 sky130_fd_sc_hd__clkbuf_1 _20308_ (.A(_04724_),
    .X(_00957_));
 sky130_fd_sc_hd__nand2_1 _20309_ (.A(_04715_),
    .B(_12214_),
    .Y(_04725_));
 sky130_fd_sc_hd__o211a_1 _20310_ (.A1(_03236_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _20311_ (.A0(_04726_),
    .A1(net2455),
    .S(_04705_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _20312_ (.A(_04727_),
    .X(_00958_));
 sky130_fd_sc_hd__nand2_1 _20313_ (.A(_04715_),
    .B(_12222_),
    .Y(_04728_));
 sky130_fd_sc_hd__o211a_1 _20314_ (.A1(_03240_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__mux2_1 _20315_ (.A0(_04729_),
    .A1(net3783),
    .S(_04705_),
    .X(_04730_));
 sky130_fd_sc_hd__clkbuf_1 _20316_ (.A(_04730_),
    .X(_00959_));
 sky130_fd_sc_hd__nand2_1 _20317_ (.A(_04715_),
    .B(_12230_),
    .Y(_04731_));
 sky130_fd_sc_hd__o211a_1 _20318_ (.A1(_03244_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_1 _20319_ (.A0(_04732_),
    .A1(net2522),
    .S(_04705_),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_1 _20320_ (.A(_04733_),
    .X(_00960_));
 sky130_fd_sc_hd__nand2_1 _20321_ (.A(_04715_),
    .B(_12238_),
    .Y(_04734_));
 sky130_fd_sc_hd__o211a_1 _20322_ (.A1(_03248_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _20323_ (.A0(_04735_),
    .A1(net2779),
    .S(_04705_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_1 _20324_ (.A(_04736_),
    .X(_00961_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_04715_),
    .B(_12246_),
    .Y(_04737_));
 sky130_fd_sc_hd__o211a_1 _20326_ (.A1(_03252_),
    .A2(_04714_),
    .B1(_04463_),
    .C1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__mux2_1 _20327_ (.A0(_04738_),
    .A1(net2154),
    .S(_04705_),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_1 _20328_ (.A(_04739_),
    .X(_00962_));
 sky130_fd_sc_hd__buf_4 _20329_ (.A(_03702_),
    .X(_04740_));
 sky130_fd_sc_hd__o211a_1 _20330_ (.A1(_03256_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04716_),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_8 _20331_ (.A(_04704_),
    .X(_04742_));
 sky130_fd_sc_hd__mux2_1 _20332_ (.A0(_04741_),
    .A1(net2749),
    .S(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_1 _20333_ (.A(_04743_),
    .X(_00963_));
 sky130_fd_sc_hd__o211a_1 _20334_ (.A1(_03261_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04719_),
    .X(_04744_));
 sky130_fd_sc_hd__mux2_1 _20335_ (.A0(_04744_),
    .A1(net3472),
    .S(_04742_),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_1 _20336_ (.A(_04745_),
    .X(_00964_));
 sky130_fd_sc_hd__o211a_1 _20337_ (.A1(_03264_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04722_),
    .X(_04746_));
 sky130_fd_sc_hd__mux2_1 _20338_ (.A0(_04746_),
    .A1(net3621),
    .S(_04742_),
    .X(_04747_));
 sky130_fd_sc_hd__clkbuf_1 _20339_ (.A(_04747_),
    .X(_00965_));
 sky130_fd_sc_hd__o211a_1 _20340_ (.A1(_03267_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04725_),
    .X(_04748_));
 sky130_fd_sc_hd__mux2_1 _20341_ (.A0(_04748_),
    .A1(net3119),
    .S(_04742_),
    .X(_04749_));
 sky130_fd_sc_hd__clkbuf_1 _20342_ (.A(_04749_),
    .X(_00966_));
 sky130_fd_sc_hd__o211a_1 _20343_ (.A1(_03270_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04728_),
    .X(_04750_));
 sky130_fd_sc_hd__mux2_1 _20344_ (.A0(_04750_),
    .A1(net3684),
    .S(_04742_),
    .X(_04751_));
 sky130_fd_sc_hd__clkbuf_1 _20345_ (.A(_04751_),
    .X(_00967_));
 sky130_fd_sc_hd__o211a_1 _20346_ (.A1(_03273_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04731_),
    .X(_04752_));
 sky130_fd_sc_hd__mux2_1 _20347_ (.A0(_04752_),
    .A1(net2815),
    .S(_04742_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_1 _20348_ (.A(_04753_),
    .X(_00968_));
 sky130_fd_sc_hd__o211a_1 _20349_ (.A1(_03276_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04734_),
    .X(_04754_));
 sky130_fd_sc_hd__mux2_1 _20350_ (.A0(_04754_),
    .A1(net3556),
    .S(_04742_),
    .X(_04755_));
 sky130_fd_sc_hd__clkbuf_1 _20351_ (.A(_04755_),
    .X(_00969_));
 sky130_fd_sc_hd__o211a_1 _20352_ (.A1(_03279_),
    .A2(_04714_),
    .B1(_04740_),
    .C1(_04737_),
    .X(_04756_));
 sky130_fd_sc_hd__mux2_1 _20353_ (.A0(_04756_),
    .A1(net3248),
    .S(_04742_),
    .X(_04757_));
 sky130_fd_sc_hd__clkbuf_1 _20354_ (.A(_04757_),
    .X(_00970_));
 sky130_fd_sc_hd__o211a_1 _20355_ (.A1(_12170_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04716_),
    .X(_04758_));
 sky130_fd_sc_hd__mux2_1 _20356_ (.A0(_04758_),
    .A1(net2324),
    .S(_04742_),
    .X(_04759_));
 sky130_fd_sc_hd__clkbuf_1 _20357_ (.A(_04759_),
    .X(_00971_));
 sky130_fd_sc_hd__o211a_1 _20358_ (.A1(_12195_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04719_),
    .X(_04760_));
 sky130_fd_sc_hd__mux2_1 _20359_ (.A0(_04760_),
    .A1(net2158),
    .S(_04742_),
    .X(_04761_));
 sky130_fd_sc_hd__clkbuf_1 _20360_ (.A(_04761_),
    .X(_00972_));
 sky130_fd_sc_hd__o211a_1 _20361_ (.A1(_12203_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04722_),
    .X(_04762_));
 sky130_fd_sc_hd__mux2_1 _20362_ (.A0(_04762_),
    .A1(net2697),
    .S(_04742_),
    .X(_04763_));
 sky130_fd_sc_hd__clkbuf_1 _20363_ (.A(_04763_),
    .X(_00973_));
 sky130_fd_sc_hd__o211a_1 _20364_ (.A1(_12211_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04725_),
    .X(_04764_));
 sky130_fd_sc_hd__mux2_1 _20365_ (.A0(_04764_),
    .A1(net2382),
    .S(_04742_),
    .X(_04765_));
 sky130_fd_sc_hd__clkbuf_1 _20366_ (.A(_04765_),
    .X(_00974_));
 sky130_fd_sc_hd__o211a_1 _20367_ (.A1(_12219_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04728_),
    .X(_04766_));
 sky130_fd_sc_hd__mux2_1 _20368_ (.A0(_04766_),
    .A1(net3760),
    .S(_04742_),
    .X(_04767_));
 sky130_fd_sc_hd__clkbuf_1 _20369_ (.A(_04767_),
    .X(_00975_));
 sky130_fd_sc_hd__o211a_1 _20370_ (.A1(_12227_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04731_),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_1 _20371_ (.A0(_04768_),
    .A1(net2908),
    .S(_04742_),
    .X(_04769_));
 sky130_fd_sc_hd__clkbuf_1 _20372_ (.A(_04769_),
    .X(_00976_));
 sky130_fd_sc_hd__o211a_1 _20373_ (.A1(_12235_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04734_),
    .X(_04770_));
 sky130_fd_sc_hd__mux2_1 _20374_ (.A0(_04770_),
    .A1(net3229),
    .S(_04742_),
    .X(_04771_));
 sky130_fd_sc_hd__clkbuf_1 _20375_ (.A(_04771_),
    .X(_00977_));
 sky130_fd_sc_hd__o211a_1 _20376_ (.A1(_12243_),
    .A2(_04715_),
    .B1(_04740_),
    .C1(_04737_),
    .X(_04772_));
 sky130_fd_sc_hd__mux2_1 _20377_ (.A0(_04772_),
    .A1(net3296),
    .S(_04742_),
    .X(_04773_));
 sky130_fd_sc_hd__clkbuf_1 _20378_ (.A(_04773_),
    .X(_00978_));
 sky130_fd_sc_hd__nand2_1 _20379_ (.A(_04702_),
    .B(_04183_),
    .Y(_04774_));
 sky130_fd_sc_hd__inv_2 _20380_ (.A(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__clkbuf_16 _20381_ (.A(_12190_),
    .X(_04776_));
 sky130_fd_sc_hd__o21ai_4 _20382_ (.A1(_04332_),
    .A2(_04775_),
    .B1(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__mux2_1 _20383_ (.A0(_04101_),
    .A1(net2663),
    .S(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__clkbuf_1 _20384_ (.A(_04778_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _20385_ (.A0(_04109_),
    .A1(net2549),
    .S(_04777_),
    .X(_04779_));
 sky130_fd_sc_hd__clkbuf_1 _20386_ (.A(_04779_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _20387_ (.A0(_04111_),
    .A1(net3471),
    .S(_04777_),
    .X(_04780_));
 sky130_fd_sc_hd__clkbuf_1 _20388_ (.A(_04780_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _20389_ (.A0(_04113_),
    .A1(net3130),
    .S(_04777_),
    .X(_04781_));
 sky130_fd_sc_hd__clkbuf_1 _20390_ (.A(_04781_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _20391_ (.A0(_04115_),
    .A1(net3044),
    .S(_04777_),
    .X(_04782_));
 sky130_fd_sc_hd__clkbuf_1 _20392_ (.A(_04782_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _20393_ (.A0(_04117_),
    .A1(net2738),
    .S(_04777_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_1 _20394_ (.A(_04783_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _20395_ (.A0(_04119_),
    .A1(net3216),
    .S(_04777_),
    .X(_04784_));
 sky130_fd_sc_hd__clkbuf_1 _20396_ (.A(_04784_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _20397_ (.A0(_04121_),
    .A1(net3186),
    .S(_04777_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_1 _20398_ (.A(_04785_),
    .X(_00986_));
 sky130_fd_sc_hd__buf_4 _20399_ (.A(_04777_),
    .X(_04786_));
 sky130_fd_sc_hd__buf_4 _20400_ (.A(_04775_),
    .X(_04787_));
 sky130_fd_sc_hd__buf_4 _20401_ (.A(_04775_),
    .X(_04788_));
 sky130_fd_sc_hd__nor2_1 _20402_ (.A(_02854_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__a211o_1 _20403_ (.A1(_02852_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__buf_4 _20404_ (.A(_04777_),
    .X(_04791_));
 sky130_fd_sc_hd__nand2_1 _20405_ (.A(_04791_),
    .B(net890),
    .Y(_04792_));
 sky130_fd_sc_hd__o21ai_1 _20406_ (.A1(_04786_),
    .A2(_04790_),
    .B1(net891),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _20407_ (.A(_02863_),
    .B(_04788_),
    .Y(_04793_));
 sky130_fd_sc_hd__a211o_1 _20408_ (.A1(_02862_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__nand2_1 _20409_ (.A(_04791_),
    .B(net1498),
    .Y(_04795_));
 sky130_fd_sc_hd__o21ai_1 _20410_ (.A1(_04786_),
    .A2(_04794_),
    .B1(net1499),
    .Y(_00988_));
 sky130_fd_sc_hd__nor2_1 _20411_ (.A(_02870_),
    .B(_04788_),
    .Y(_04796_));
 sky130_fd_sc_hd__a211o_1 _20412_ (.A1(_02869_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__nand2_1 _20413_ (.A(_04791_),
    .B(net682),
    .Y(_04798_));
 sky130_fd_sc_hd__o21ai_1 _20414_ (.A1(_04786_),
    .A2(_04797_),
    .B1(net683),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _20415_ (.A(_02877_),
    .B(_04788_),
    .Y(_04799_));
 sky130_fd_sc_hd__a211o_1 _20416_ (.A1(_02876_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_1 _20417_ (.A(_04791_),
    .B(net1106),
    .Y(_04801_));
 sky130_fd_sc_hd__o21ai_1 _20418_ (.A1(_04786_),
    .A2(_04800_),
    .B1(net1107),
    .Y(_00990_));
 sky130_fd_sc_hd__nor2_1 _20419_ (.A(_02884_),
    .B(_04788_),
    .Y(_04802_));
 sky130_fd_sc_hd__a211o_1 _20420_ (.A1(_02883_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__nand2_1 _20421_ (.A(_04791_),
    .B(net984),
    .Y(_04804_));
 sky130_fd_sc_hd__o21ai_1 _20422_ (.A1(_04786_),
    .A2(_04803_),
    .B1(net985),
    .Y(_00991_));
 sky130_fd_sc_hd__nor2_1 _20423_ (.A(_02891_),
    .B(_04788_),
    .Y(_04805_));
 sky130_fd_sc_hd__a211o_1 _20424_ (.A1(_02890_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__nand2_1 _20425_ (.A(_04791_),
    .B(net1208),
    .Y(_04807_));
 sky130_fd_sc_hd__o21ai_1 _20426_ (.A1(_04786_),
    .A2(_04806_),
    .B1(net1209),
    .Y(_00992_));
 sky130_fd_sc_hd__nor2_1 _20427_ (.A(_02898_),
    .B(_04788_),
    .Y(_04808_));
 sky130_fd_sc_hd__a211o_1 _20428_ (.A1(_02897_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__nand2_1 _20429_ (.A(_04791_),
    .B(net806),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ai_1 _20430_ (.A1(_04786_),
    .A2(_04809_),
    .B1(net807),
    .Y(_00993_));
 sky130_fd_sc_hd__nor2_1 _20431_ (.A(_02905_),
    .B(_04788_),
    .Y(_04811_));
 sky130_fd_sc_hd__a211o_1 _20432_ (.A1(_02904_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__nand2_1 _20433_ (.A(_04791_),
    .B(net1238),
    .Y(_04813_));
 sky130_fd_sc_hd__o21ai_1 _20434_ (.A1(_04786_),
    .A2(_04812_),
    .B1(net1239),
    .Y(_00994_));
 sky130_fd_sc_hd__buf_4 _20435_ (.A(_04777_),
    .X(_04814_));
 sky130_fd_sc_hd__a211o_1 _20436_ (.A1(_02912_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04789_),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_1 _20437_ (.A(_04791_),
    .B(net1390),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ai_1 _20438_ (.A1(_04814_),
    .A2(_04815_),
    .B1(net1391),
    .Y(_00995_));
 sky130_fd_sc_hd__a211o_1 _20439_ (.A1(_02917_),
    .A2(_04787_),
    .B1(_04689_),
    .C1(_04793_),
    .X(_04817_));
 sky130_fd_sc_hd__nand2_1 _20440_ (.A(_04791_),
    .B(net1610),
    .Y(_04818_));
 sky130_fd_sc_hd__o21ai_1 _20441_ (.A1(_04814_),
    .A2(_04817_),
    .B1(net1611),
    .Y(_00996_));
 sky130_fd_sc_hd__buf_4 _20442_ (.A(_04598_),
    .X(_04819_));
 sky130_fd_sc_hd__a211o_1 _20443_ (.A1(_02922_),
    .A2(_04787_),
    .B1(_04819_),
    .C1(_04796_),
    .X(_04820_));
 sky130_fd_sc_hd__nand2_1 _20444_ (.A(_04791_),
    .B(net1848),
    .Y(_04821_));
 sky130_fd_sc_hd__o21ai_1 _20445_ (.A1(_04814_),
    .A2(_04820_),
    .B1(net1849),
    .Y(_00997_));
 sky130_fd_sc_hd__a211o_1 _20446_ (.A1(_02928_),
    .A2(_04787_),
    .B1(_04819_),
    .C1(_04799_),
    .X(_04822_));
 sky130_fd_sc_hd__nand2_1 _20447_ (.A(_04791_),
    .B(net1288),
    .Y(_04823_));
 sky130_fd_sc_hd__o21ai_1 _20448_ (.A1(_04814_),
    .A2(_04822_),
    .B1(net1289),
    .Y(_00998_));
 sky130_fd_sc_hd__a211o_1 _20449_ (.A1(_02933_),
    .A2(_04787_),
    .B1(_04819_),
    .C1(_04802_),
    .X(_04824_));
 sky130_fd_sc_hd__nand2_1 _20450_ (.A(_04791_),
    .B(net1764),
    .Y(_04825_));
 sky130_fd_sc_hd__o21ai_1 _20451_ (.A1(_04814_),
    .A2(_04824_),
    .B1(net1765),
    .Y(_00999_));
 sky130_fd_sc_hd__a211o_1 _20452_ (.A1(_02938_),
    .A2(_04787_),
    .B1(_04819_),
    .C1(_04805_),
    .X(_04826_));
 sky130_fd_sc_hd__nand2_1 _20453_ (.A(_04791_),
    .B(net1744),
    .Y(_04827_));
 sky130_fd_sc_hd__o21ai_1 _20454_ (.A1(_04814_),
    .A2(_04826_),
    .B1(net1745),
    .Y(_01000_));
 sky130_fd_sc_hd__a211o_1 _20455_ (.A1(_02943_),
    .A2(_04787_),
    .B1(_04819_),
    .C1(_04808_),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_1 _20456_ (.A(_04791_),
    .B(net1712),
    .Y(_04829_));
 sky130_fd_sc_hd__o21ai_1 _20457_ (.A1(_04814_),
    .A2(_04828_),
    .B1(net1713),
    .Y(_01001_));
 sky130_fd_sc_hd__a211o_1 _20458_ (.A1(_02948_),
    .A2(_04787_),
    .B1(_04819_),
    .C1(_04811_),
    .X(_04830_));
 sky130_fd_sc_hd__nand2_1 _20459_ (.A(_04791_),
    .B(net1620),
    .Y(_04831_));
 sky130_fd_sc_hd__o21ai_1 _20460_ (.A1(_04814_),
    .A2(_04830_),
    .B1(net1621),
    .Y(_01002_));
 sky130_fd_sc_hd__a211o_1 _20461_ (.A1(_02952_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04789_),
    .X(_04832_));
 sky130_fd_sc_hd__nand2_1 _20462_ (.A(_04786_),
    .B(net556),
    .Y(_04833_));
 sky130_fd_sc_hd__o21ai_1 _20463_ (.A1(_04814_),
    .A2(_04832_),
    .B1(net557),
    .Y(_01003_));
 sky130_fd_sc_hd__a211o_1 _20464_ (.A1(_02956_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04793_),
    .X(_04834_));
 sky130_fd_sc_hd__nand2_1 _20465_ (.A(_04786_),
    .B(net1086),
    .Y(_04835_));
 sky130_fd_sc_hd__o21ai_1 _20466_ (.A1(_04814_),
    .A2(_04834_),
    .B1(net1087),
    .Y(_01004_));
 sky130_fd_sc_hd__a211o_1 _20467_ (.A1(_02960_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04796_),
    .X(_04836_));
 sky130_fd_sc_hd__nand2_1 _20468_ (.A(_04786_),
    .B(net1078),
    .Y(_04837_));
 sky130_fd_sc_hd__o21ai_1 _20469_ (.A1(_04814_),
    .A2(_04836_),
    .B1(net1079),
    .Y(_01005_));
 sky130_fd_sc_hd__a211o_1 _20470_ (.A1(_02964_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04799_),
    .X(_04838_));
 sky130_fd_sc_hd__nand2_1 _20471_ (.A(_04786_),
    .B(net1334),
    .Y(_04839_));
 sky130_fd_sc_hd__o21ai_1 _20472_ (.A1(_04814_),
    .A2(_04838_),
    .B1(net1335),
    .Y(_01006_));
 sky130_fd_sc_hd__a211o_1 _20473_ (.A1(_02968_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04802_),
    .X(_04840_));
 sky130_fd_sc_hd__nand2_1 _20474_ (.A(_04786_),
    .B(net728),
    .Y(_04841_));
 sky130_fd_sc_hd__o21ai_1 _20475_ (.A1(_04814_),
    .A2(_04840_),
    .B1(net729),
    .Y(_01007_));
 sky130_fd_sc_hd__a211o_1 _20476_ (.A1(_02972_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04805_),
    .X(_04842_));
 sky130_fd_sc_hd__nand2_1 _20477_ (.A(_04786_),
    .B(net1372),
    .Y(_04843_));
 sky130_fd_sc_hd__o21ai_1 _20478_ (.A1(_04814_),
    .A2(_04842_),
    .B1(net1373),
    .Y(_01008_));
 sky130_fd_sc_hd__a211o_1 _20479_ (.A1(_02976_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04808_),
    .X(_04844_));
 sky130_fd_sc_hd__nand2_1 _20480_ (.A(_04786_),
    .B(net1240),
    .Y(_04845_));
 sky130_fd_sc_hd__o21ai_1 _20481_ (.A1(_04814_),
    .A2(_04844_),
    .B1(net1241),
    .Y(_01009_));
 sky130_fd_sc_hd__a211o_1 _20482_ (.A1(_02980_),
    .A2(_04788_),
    .B1(_04819_),
    .C1(_04811_),
    .X(_04846_));
 sky130_fd_sc_hd__nand2_1 _20483_ (.A(_04786_),
    .B(net942),
    .Y(_04847_));
 sky130_fd_sc_hd__o21ai_1 _20484_ (.A1(_04814_),
    .A2(_04846_),
    .B1(net943),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _20485_ (.A(_04702_),
    .B(_04257_),
    .Y(_04848_));
 sky130_fd_sc_hd__inv_2 _20486_ (.A(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__o21ai_4 _20487_ (.A1(_04332_),
    .A2(_04849_),
    .B1(_04776_),
    .Y(_04850_));
 sky130_fd_sc_hd__mux2_1 _20488_ (.A0(_04101_),
    .A1(net2437),
    .S(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_1 _20489_ (.A(_04851_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _20490_ (.A0(_04109_),
    .A1(net2031),
    .S(_04850_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _20491_ (.A(_04852_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _20492_ (.A0(_04111_),
    .A1(net2195),
    .S(_04850_),
    .X(_04853_));
 sky130_fd_sc_hd__clkbuf_1 _20493_ (.A(_04853_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _20494_ (.A0(_04113_),
    .A1(net2137),
    .S(_04850_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_1 _20495_ (.A(_04854_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _20496_ (.A0(_04115_),
    .A1(net2634),
    .S(_04850_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_1 _20497_ (.A(_04855_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _20498_ (.A0(_04117_),
    .A1(net2162),
    .S(_04850_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_1 _20499_ (.A(_04856_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _20500_ (.A0(_04119_),
    .A1(net2099),
    .S(_04850_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _20501_ (.A(_04857_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _20502_ (.A0(_04121_),
    .A1(net2138),
    .S(_04850_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_1 _20503_ (.A(_04858_),
    .X(_01018_));
 sky130_fd_sc_hd__buf_4 _20504_ (.A(_04850_),
    .X(_04859_));
 sky130_fd_sc_hd__buf_4 _20505_ (.A(_04849_),
    .X(_04860_));
 sky130_fd_sc_hd__buf_4 _20506_ (.A(_04849_),
    .X(_04861_));
 sky130_fd_sc_hd__nor2_1 _20507_ (.A(_02854_),
    .B(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__a211o_1 _20508_ (.A1(_02852_),
    .A2(_04860_),
    .B1(_04819_),
    .C1(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__buf_4 _20509_ (.A(_04850_),
    .X(_04864_));
 sky130_fd_sc_hd__nand2_1 _20510_ (.A(_04864_),
    .B(net788),
    .Y(_04865_));
 sky130_fd_sc_hd__o21ai_1 _20511_ (.A1(_04859_),
    .A2(_04863_),
    .B1(net789),
    .Y(_01019_));
 sky130_fd_sc_hd__nor2_1 _20512_ (.A(_02863_),
    .B(_04861_),
    .Y(_04866_));
 sky130_fd_sc_hd__a211o_1 _20513_ (.A1(_02862_),
    .A2(_04860_),
    .B1(_04819_),
    .C1(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_1 _20514_ (.A(_04864_),
    .B(net418),
    .Y(_04868_));
 sky130_fd_sc_hd__o21ai_1 _20515_ (.A1(_04859_),
    .A2(_04867_),
    .B1(net419),
    .Y(_01020_));
 sky130_fd_sc_hd__buf_4 _20516_ (.A(_04598_),
    .X(_04869_));
 sky130_fd_sc_hd__nor2_1 _20517_ (.A(_02870_),
    .B(_04861_),
    .Y(_04870_));
 sky130_fd_sc_hd__a211o_1 _20518_ (.A1(_02869_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__nand2_1 _20519_ (.A(_04864_),
    .B(net404),
    .Y(_04872_));
 sky130_fd_sc_hd__o21ai_1 _20520_ (.A1(_04859_),
    .A2(_04871_),
    .B1(net405),
    .Y(_01021_));
 sky130_fd_sc_hd__nor2_1 _20521_ (.A(_02877_),
    .B(_04861_),
    .Y(_04873_));
 sky130_fd_sc_hd__a211o_1 _20522_ (.A1(_02876_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _20523_ (.A(_04864_),
    .B(net510),
    .Y(_04875_));
 sky130_fd_sc_hd__o21ai_1 _20524_ (.A1(_04859_),
    .A2(_04874_),
    .B1(net511),
    .Y(_01022_));
 sky130_fd_sc_hd__nor2_1 _20525_ (.A(_02884_),
    .B(_04861_),
    .Y(_04876_));
 sky130_fd_sc_hd__a211o_1 _20526_ (.A1(_02883_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__nand2_1 _20527_ (.A(_04864_),
    .B(net524),
    .Y(_04878_));
 sky130_fd_sc_hd__o21ai_1 _20528_ (.A1(_04859_),
    .A2(_04877_),
    .B1(net525),
    .Y(_01023_));
 sky130_fd_sc_hd__nor2_1 _20529_ (.A(_02891_),
    .B(_04861_),
    .Y(_04879_));
 sky130_fd_sc_hd__a211o_1 _20530_ (.A1(_02890_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__nand2_1 _20531_ (.A(_04864_),
    .B(net960),
    .Y(_04881_));
 sky130_fd_sc_hd__o21ai_1 _20532_ (.A1(_04859_),
    .A2(_04880_),
    .B1(net961),
    .Y(_01024_));
 sky130_fd_sc_hd__nor2_1 _20533_ (.A(_02898_),
    .B(_04861_),
    .Y(_04882_));
 sky130_fd_sc_hd__a211o_1 _20534_ (.A1(_02897_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__nand2_1 _20535_ (.A(_04864_),
    .B(net390),
    .Y(_04884_));
 sky130_fd_sc_hd__o21ai_1 _20536_ (.A1(_04859_),
    .A2(_04883_),
    .B1(net391),
    .Y(_01025_));
 sky130_fd_sc_hd__nor2_1 _20537_ (.A(_02905_),
    .B(_04861_),
    .Y(_04885_));
 sky130_fd_sc_hd__a211o_1 _20538_ (.A1(_02904_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__nand2_1 _20539_ (.A(_04864_),
    .B(net494),
    .Y(_04887_));
 sky130_fd_sc_hd__o21ai_1 _20540_ (.A1(_04859_),
    .A2(_04886_),
    .B1(net495),
    .Y(_01026_));
 sky130_fd_sc_hd__buf_4 _20541_ (.A(_04850_),
    .X(_04888_));
 sky130_fd_sc_hd__a211o_1 _20542_ (.A1(_02912_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04862_),
    .X(_04889_));
 sky130_fd_sc_hd__nand2_1 _20543_ (.A(_04864_),
    .B(net542),
    .Y(_04890_));
 sky130_fd_sc_hd__o21ai_1 _20544_ (.A1(_04888_),
    .A2(_04889_),
    .B1(net543),
    .Y(_01027_));
 sky130_fd_sc_hd__a211o_1 _20545_ (.A1(_02917_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04866_),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_1 _20546_ (.A(_04864_),
    .B(net426),
    .Y(_04892_));
 sky130_fd_sc_hd__o21ai_1 _20547_ (.A1(_04888_),
    .A2(_04891_),
    .B1(net427),
    .Y(_01028_));
 sky130_fd_sc_hd__a211o_1 _20548_ (.A1(_02922_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04870_),
    .X(_04893_));
 sky130_fd_sc_hd__nand2_1 _20549_ (.A(_04864_),
    .B(net794),
    .Y(_04894_));
 sky130_fd_sc_hd__o21ai_1 _20550_ (.A1(_04888_),
    .A2(_04893_),
    .B1(net795),
    .Y(_01029_));
 sky130_fd_sc_hd__a211o_1 _20551_ (.A1(_02928_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04873_),
    .X(_04895_));
 sky130_fd_sc_hd__nand2_1 _20552_ (.A(_04864_),
    .B(net504),
    .Y(_04896_));
 sky130_fd_sc_hd__o21ai_1 _20553_ (.A1(_04888_),
    .A2(_04895_),
    .B1(net505),
    .Y(_01030_));
 sky130_fd_sc_hd__a211o_1 _20554_ (.A1(_02933_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04876_),
    .X(_04897_));
 sky130_fd_sc_hd__nand2_1 _20555_ (.A(_04864_),
    .B(net762),
    .Y(_04898_));
 sky130_fd_sc_hd__o21ai_1 _20556_ (.A1(_04888_),
    .A2(_04897_),
    .B1(net763),
    .Y(_01031_));
 sky130_fd_sc_hd__a211o_1 _20557_ (.A1(_02938_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04879_),
    .X(_04899_));
 sky130_fd_sc_hd__nand2_1 _20558_ (.A(_04864_),
    .B(net526),
    .Y(_04900_));
 sky130_fd_sc_hd__o21ai_1 _20559_ (.A1(_04888_),
    .A2(_04899_),
    .B1(net527),
    .Y(_01032_));
 sky130_fd_sc_hd__a211o_1 _20560_ (.A1(_02943_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04882_),
    .X(_04901_));
 sky130_fd_sc_hd__nand2_1 _20561_ (.A(_04864_),
    .B(net444),
    .Y(_04902_));
 sky130_fd_sc_hd__o21ai_1 _20562_ (.A1(_04888_),
    .A2(_04901_),
    .B1(net445),
    .Y(_01033_));
 sky130_fd_sc_hd__a211o_1 _20563_ (.A1(_02948_),
    .A2(_04860_),
    .B1(_04869_),
    .C1(_04885_),
    .X(_04903_));
 sky130_fd_sc_hd__nand2_1 _20564_ (.A(_04864_),
    .B(net460),
    .Y(_04904_));
 sky130_fd_sc_hd__o21ai_1 _20565_ (.A1(_04888_),
    .A2(_04903_),
    .B1(net461),
    .Y(_01034_));
 sky130_fd_sc_hd__a211o_1 _20566_ (.A1(_02952_),
    .A2(_04861_),
    .B1(_04869_),
    .C1(_04862_),
    .X(_04905_));
 sky130_fd_sc_hd__nand2_1 _20567_ (.A(_04859_),
    .B(net674),
    .Y(_04906_));
 sky130_fd_sc_hd__o21ai_1 _20568_ (.A1(_04888_),
    .A2(_04905_),
    .B1(net675),
    .Y(_01035_));
 sky130_fd_sc_hd__a211o_1 _20569_ (.A1(_02956_),
    .A2(_04861_),
    .B1(_04869_),
    .C1(_04866_),
    .X(_04907_));
 sky130_fd_sc_hd__nand2_1 _20570_ (.A(_04859_),
    .B(net506),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ai_1 _20571_ (.A1(_04888_),
    .A2(_04907_),
    .B1(net507),
    .Y(_01036_));
 sky130_fd_sc_hd__clkbuf_8 _20572_ (.A(_04598_),
    .X(_04909_));
 sky130_fd_sc_hd__a211o_1 _20573_ (.A1(_02960_),
    .A2(_04861_),
    .B1(_04909_),
    .C1(_04870_),
    .X(_04910_));
 sky130_fd_sc_hd__nand2_1 _20574_ (.A(_04859_),
    .B(net602),
    .Y(_04911_));
 sky130_fd_sc_hd__o21ai_1 _20575_ (.A1(_04888_),
    .A2(_04910_),
    .B1(net603),
    .Y(_01037_));
 sky130_fd_sc_hd__a211o_1 _20576_ (.A1(_02964_),
    .A2(_04861_),
    .B1(_04909_),
    .C1(_04873_),
    .X(_04912_));
 sky130_fd_sc_hd__nand2_1 _20577_ (.A(_04859_),
    .B(net438),
    .Y(_04913_));
 sky130_fd_sc_hd__o21ai_1 _20578_ (.A1(_04888_),
    .A2(_04912_),
    .B1(net439),
    .Y(_01038_));
 sky130_fd_sc_hd__a211o_1 _20579_ (.A1(_02968_),
    .A2(_04861_),
    .B1(_04909_),
    .C1(_04876_),
    .X(_04914_));
 sky130_fd_sc_hd__nand2_1 _20580_ (.A(_04859_),
    .B(net592),
    .Y(_04915_));
 sky130_fd_sc_hd__o21ai_1 _20581_ (.A1(_04888_),
    .A2(_04914_),
    .B1(net593),
    .Y(_01039_));
 sky130_fd_sc_hd__a211o_1 _20582_ (.A1(_02972_),
    .A2(_04861_),
    .B1(_04909_),
    .C1(_04879_),
    .X(_04916_));
 sky130_fd_sc_hd__nand2_1 _20583_ (.A(_04859_),
    .B(net1120),
    .Y(_04917_));
 sky130_fd_sc_hd__o21ai_1 _20584_ (.A1(_04888_),
    .A2(_04916_),
    .B1(net1121),
    .Y(_01040_));
 sky130_fd_sc_hd__a211o_1 _20585_ (.A1(_02976_),
    .A2(_04861_),
    .B1(_04909_),
    .C1(_04882_),
    .X(_04918_));
 sky130_fd_sc_hd__nand2_1 _20586_ (.A(_04859_),
    .B(net450),
    .Y(_04919_));
 sky130_fd_sc_hd__o21ai_1 _20587_ (.A1(_04888_),
    .A2(_04918_),
    .B1(net451),
    .Y(_01041_));
 sky130_fd_sc_hd__a211o_1 _20588_ (.A1(_02980_),
    .A2(_04861_),
    .B1(_04909_),
    .C1(_04885_),
    .X(_04920_));
 sky130_fd_sc_hd__nand2_1 _20589_ (.A(_04859_),
    .B(net568),
    .Y(_04921_));
 sky130_fd_sc_hd__o21ai_1 _20590_ (.A1(_04888_),
    .A2(_04920_),
    .B1(net569),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _20591_ (.A(_04702_),
    .B(_04333_),
    .Y(_04922_));
 sky130_fd_sc_hd__inv_2 _20592_ (.A(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__o21ai_4 _20593_ (.A1(_04332_),
    .A2(_04923_),
    .B1(_04776_),
    .Y(_04924_));
 sky130_fd_sc_hd__mux2_1 _20594_ (.A0(_04101_),
    .A1(net2794),
    .S(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__clkbuf_1 _20595_ (.A(_04925_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _20596_ (.A0(_04109_),
    .A1(net3627),
    .S(_04924_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _20597_ (.A(_04926_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _20598_ (.A0(_04111_),
    .A1(net2685),
    .S(_04924_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_1 _20599_ (.A(_04927_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _20600_ (.A0(_04113_),
    .A1(net3811),
    .S(_04924_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_1 _20601_ (.A(_04928_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _20602_ (.A0(_04115_),
    .A1(net3075),
    .S(_04924_),
    .X(_04929_));
 sky130_fd_sc_hd__clkbuf_1 _20603_ (.A(_04929_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _20604_ (.A0(_04117_),
    .A1(net2996),
    .S(_04924_),
    .X(_04930_));
 sky130_fd_sc_hd__clkbuf_1 _20605_ (.A(_04930_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _20606_ (.A0(_04119_),
    .A1(net3210),
    .S(_04924_),
    .X(_04931_));
 sky130_fd_sc_hd__clkbuf_1 _20607_ (.A(_04931_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _20608_ (.A0(_04121_),
    .A1(net2581),
    .S(_04924_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_1 _20609_ (.A(_04932_),
    .X(_01050_));
 sky130_fd_sc_hd__buf_4 _20610_ (.A(_04924_),
    .X(_04933_));
 sky130_fd_sc_hd__buf_4 _20611_ (.A(_04923_),
    .X(_04934_));
 sky130_fd_sc_hd__buf_4 _20612_ (.A(_04923_),
    .X(_04935_));
 sky130_fd_sc_hd__nor2_1 _20613_ (.A(_02854_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__a211o_1 _20614_ (.A1(_02852_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__buf_4 _20615_ (.A(_04924_),
    .X(_04938_));
 sky130_fd_sc_hd__nand2_1 _20616_ (.A(_04938_),
    .B(net1038),
    .Y(_04939_));
 sky130_fd_sc_hd__o21ai_1 _20617_ (.A1(_04933_),
    .A2(_04937_),
    .B1(net1039),
    .Y(_01051_));
 sky130_fd_sc_hd__nor2_1 _20618_ (.A(_02863_),
    .B(_04935_),
    .Y(_04940_));
 sky130_fd_sc_hd__a211o_1 _20619_ (.A1(_02862_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _20620_ (.A(_04938_),
    .B(net580),
    .Y(_04942_));
 sky130_fd_sc_hd__o21ai_1 _20621_ (.A1(_04933_),
    .A2(_04941_),
    .B1(net581),
    .Y(_01052_));
 sky130_fd_sc_hd__nor2_1 _20622_ (.A(_02870_),
    .B(_04935_),
    .Y(_04943_));
 sky130_fd_sc_hd__a211o_1 _20623_ (.A1(_02869_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__nand2_1 _20624_ (.A(_04938_),
    .B(net1446),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ai_1 _20625_ (.A1(_04933_),
    .A2(_04944_),
    .B1(net1447),
    .Y(_01053_));
 sky130_fd_sc_hd__nor2_1 _20626_ (.A(_02877_),
    .B(_04935_),
    .Y(_04946_));
 sky130_fd_sc_hd__a211o_1 _20627_ (.A1(_02876_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__nand2_1 _20628_ (.A(_04938_),
    .B(net1122),
    .Y(_04948_));
 sky130_fd_sc_hd__o21ai_1 _20629_ (.A1(_04933_),
    .A2(_04947_),
    .B1(net1123),
    .Y(_01054_));
 sky130_fd_sc_hd__nor2_1 _20630_ (.A(_02884_),
    .B(_04935_),
    .Y(_04949_));
 sky130_fd_sc_hd__a211o_1 _20631_ (.A1(_02883_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__nand2_1 _20632_ (.A(_04938_),
    .B(net586),
    .Y(_04951_));
 sky130_fd_sc_hd__o21ai_1 _20633_ (.A1(_04933_),
    .A2(_04950_),
    .B1(net587),
    .Y(_01055_));
 sky130_fd_sc_hd__nor2_1 _20634_ (.A(_02891_),
    .B(_04935_),
    .Y(_04952_));
 sky130_fd_sc_hd__a211o_1 _20635_ (.A1(_02890_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__nand2_1 _20636_ (.A(_04938_),
    .B(net990),
    .Y(_04954_));
 sky130_fd_sc_hd__o21ai_1 _20637_ (.A1(_04933_),
    .A2(_04953_),
    .B1(net991),
    .Y(_01056_));
 sky130_fd_sc_hd__nor2_1 _20638_ (.A(_02898_),
    .B(_04935_),
    .Y(_04955_));
 sky130_fd_sc_hd__a211o_1 _20639_ (.A1(_02897_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__nand2_1 _20640_ (.A(_04938_),
    .B(net964),
    .Y(_04957_));
 sky130_fd_sc_hd__o21ai_1 _20641_ (.A1(_04933_),
    .A2(_04956_),
    .B1(net965),
    .Y(_01057_));
 sky130_fd_sc_hd__nor2_1 _20642_ (.A(_02905_),
    .B(_04935_),
    .Y(_04958_));
 sky130_fd_sc_hd__a211o_1 _20643_ (.A1(_02904_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__nand2_1 _20644_ (.A(_04938_),
    .B(net600),
    .Y(_04960_));
 sky130_fd_sc_hd__o21ai_1 _20645_ (.A1(_04933_),
    .A2(_04959_),
    .B1(net601),
    .Y(_01058_));
 sky130_fd_sc_hd__buf_4 _20646_ (.A(_04924_),
    .X(_04961_));
 sky130_fd_sc_hd__a211o_1 _20647_ (.A1(_02912_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04936_),
    .X(_04962_));
 sky130_fd_sc_hd__nand2_1 _20648_ (.A(_04938_),
    .B(net1210),
    .Y(_04963_));
 sky130_fd_sc_hd__o21ai_1 _20649_ (.A1(_04961_),
    .A2(_04962_),
    .B1(net1211),
    .Y(_01059_));
 sky130_fd_sc_hd__a211o_1 _20650_ (.A1(_02917_),
    .A2(_04934_),
    .B1(_04909_),
    .C1(_04940_),
    .X(_04964_));
 sky130_fd_sc_hd__nand2_1 _20651_ (.A(_04938_),
    .B(net1658),
    .Y(_04965_));
 sky130_fd_sc_hd__o21ai_1 _20652_ (.A1(_04961_),
    .A2(_04964_),
    .B1(net1659),
    .Y(_01060_));
 sky130_fd_sc_hd__clkbuf_8 _20653_ (.A(_04598_),
    .X(_04966_));
 sky130_fd_sc_hd__a211o_1 _20654_ (.A1(_02922_),
    .A2(_04934_),
    .B1(_04966_),
    .C1(_04943_),
    .X(_04967_));
 sky130_fd_sc_hd__nand2_1 _20655_ (.A(_04938_),
    .B(net1252),
    .Y(_04968_));
 sky130_fd_sc_hd__o21ai_1 _20656_ (.A1(_04961_),
    .A2(_04967_),
    .B1(net1253),
    .Y(_01061_));
 sky130_fd_sc_hd__a211o_1 _20657_ (.A1(_02928_),
    .A2(_04934_),
    .B1(_04966_),
    .C1(_04946_),
    .X(_04969_));
 sky130_fd_sc_hd__nand2_1 _20658_ (.A(_04938_),
    .B(net1382),
    .Y(_04970_));
 sky130_fd_sc_hd__o21ai_1 _20659_ (.A1(_04961_),
    .A2(_04969_),
    .B1(net1383),
    .Y(_01062_));
 sky130_fd_sc_hd__a211o_1 _20660_ (.A1(_02933_),
    .A2(_04934_),
    .B1(_04966_),
    .C1(_04949_),
    .X(_04971_));
 sky130_fd_sc_hd__nand2_1 _20661_ (.A(_04938_),
    .B(net1236),
    .Y(_04972_));
 sky130_fd_sc_hd__o21ai_1 _20662_ (.A1(_04961_),
    .A2(_04971_),
    .B1(net1237),
    .Y(_01063_));
 sky130_fd_sc_hd__a211o_1 _20663_ (.A1(_02938_),
    .A2(_04934_),
    .B1(_04966_),
    .C1(_04952_),
    .X(_04973_));
 sky130_fd_sc_hd__nand2_1 _20664_ (.A(_04938_),
    .B(net666),
    .Y(_04974_));
 sky130_fd_sc_hd__o21ai_1 _20665_ (.A1(_04961_),
    .A2(_04973_),
    .B1(net667),
    .Y(_01064_));
 sky130_fd_sc_hd__a211o_1 _20666_ (.A1(_02943_),
    .A2(_04934_),
    .B1(_04966_),
    .C1(_04955_),
    .X(_04975_));
 sky130_fd_sc_hd__nand2_1 _20667_ (.A(_04938_),
    .B(net1434),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ai_1 _20668_ (.A1(_04961_),
    .A2(_04975_),
    .B1(net1435),
    .Y(_01065_));
 sky130_fd_sc_hd__a211o_1 _20669_ (.A1(_02948_),
    .A2(_04934_),
    .B1(_04966_),
    .C1(_04958_),
    .X(_04977_));
 sky130_fd_sc_hd__nand2_1 _20670_ (.A(_04938_),
    .B(net1282),
    .Y(_04978_));
 sky130_fd_sc_hd__o21ai_1 _20671_ (.A1(_04961_),
    .A2(_04977_),
    .B1(net1283),
    .Y(_01066_));
 sky130_fd_sc_hd__a211o_1 _20672_ (.A1(_02952_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04936_),
    .X(_04979_));
 sky130_fd_sc_hd__nand2_1 _20673_ (.A(_04933_),
    .B(net870),
    .Y(_04980_));
 sky130_fd_sc_hd__o21ai_1 _20674_ (.A1(_04961_),
    .A2(_04979_),
    .B1(net871),
    .Y(_01067_));
 sky130_fd_sc_hd__a211o_1 _20675_ (.A1(_02956_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04940_),
    .X(_04981_));
 sky130_fd_sc_hd__nand2_1 _20676_ (.A(_04933_),
    .B(net570),
    .Y(_04982_));
 sky130_fd_sc_hd__o21ai_1 _20677_ (.A1(_04961_),
    .A2(_04981_),
    .B1(net571),
    .Y(_01068_));
 sky130_fd_sc_hd__a211o_1 _20678_ (.A1(_02960_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04943_),
    .X(_04983_));
 sky130_fd_sc_hd__nand2_1 _20679_ (.A(_04933_),
    .B(net1284),
    .Y(_04984_));
 sky130_fd_sc_hd__o21ai_1 _20680_ (.A1(_04961_),
    .A2(_04983_),
    .B1(net1285),
    .Y(_01069_));
 sky130_fd_sc_hd__a211o_1 _20681_ (.A1(_02964_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04946_),
    .X(_04985_));
 sky130_fd_sc_hd__nand2_1 _20682_ (.A(_04933_),
    .B(net854),
    .Y(_04986_));
 sky130_fd_sc_hd__o21ai_1 _20683_ (.A1(_04961_),
    .A2(_04985_),
    .B1(net855),
    .Y(_01070_));
 sky130_fd_sc_hd__a211o_1 _20684_ (.A1(_02968_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04949_),
    .X(_04987_));
 sky130_fd_sc_hd__nand2_1 _20685_ (.A(_04933_),
    .B(net1728),
    .Y(_04988_));
 sky130_fd_sc_hd__o21ai_1 _20686_ (.A1(_04961_),
    .A2(_04987_),
    .B1(net1729),
    .Y(_01071_));
 sky130_fd_sc_hd__a211o_1 _20687_ (.A1(_02972_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04952_),
    .X(_04989_));
 sky130_fd_sc_hd__nand2_1 _20688_ (.A(_04933_),
    .B(net1594),
    .Y(_04990_));
 sky130_fd_sc_hd__o21ai_1 _20689_ (.A1(_04961_),
    .A2(_04989_),
    .B1(net1595),
    .Y(_01072_));
 sky130_fd_sc_hd__a211o_1 _20690_ (.A1(_02976_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04955_),
    .X(_04991_));
 sky130_fd_sc_hd__nand2_1 _20691_ (.A(_04933_),
    .B(net1672),
    .Y(_04992_));
 sky130_fd_sc_hd__o21ai_1 _20692_ (.A1(_04961_),
    .A2(_04991_),
    .B1(net1673),
    .Y(_01073_));
 sky130_fd_sc_hd__a211o_1 _20693_ (.A1(_02980_),
    .A2(_04935_),
    .B1(_04966_),
    .C1(_04958_),
    .X(_04993_));
 sky130_fd_sc_hd__nand2_1 _20694_ (.A(_04933_),
    .B(net760),
    .Y(_04994_));
 sky130_fd_sc_hd__o21ai_1 _20695_ (.A1(_04961_),
    .A2(_04993_),
    .B1(net761),
    .Y(_01074_));
 sky130_fd_sc_hd__and3_4 _20696_ (.A(_12173_),
    .B(_04102_),
    .C(\line_cache_idx[6] ),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_1 _20697_ (.A(_04995_),
    .B(_04104_),
    .Y(_04996_));
 sky130_fd_sc_hd__a21bo_1 _20698_ (.A1(_04996_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_04997_));
 sky130_fd_sc_hd__clkbuf_8 _20699_ (.A(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _20700_ (.A0(_04101_),
    .A1(net3110),
    .S(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__clkbuf_1 _20701_ (.A(_04999_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _20702_ (.A0(_04109_),
    .A1(net3300),
    .S(_04998_),
    .X(_05000_));
 sky130_fd_sc_hd__clkbuf_1 _20703_ (.A(_05000_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _20704_ (.A0(_04111_),
    .A1(net2864),
    .S(_04998_),
    .X(_05001_));
 sky130_fd_sc_hd__clkbuf_1 _20705_ (.A(_05001_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _20706_ (.A0(_04113_),
    .A1(net3418),
    .S(_04998_),
    .X(_05002_));
 sky130_fd_sc_hd__clkbuf_1 _20707_ (.A(_05002_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _20708_ (.A0(_04115_),
    .A1(net3196),
    .S(_04998_),
    .X(_05003_));
 sky130_fd_sc_hd__clkbuf_1 _20709_ (.A(_05003_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _20710_ (.A0(_04117_),
    .A1(net3462),
    .S(_04998_),
    .X(_05004_));
 sky130_fd_sc_hd__clkbuf_1 _20711_ (.A(_05004_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _20712_ (.A0(_04119_),
    .A1(net3436),
    .S(_04998_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_1 _20713_ (.A(_05005_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _20714_ (.A0(_04121_),
    .A1(net3098),
    .S(_04998_),
    .X(_05006_));
 sky130_fd_sc_hd__clkbuf_1 _20715_ (.A(_05006_),
    .X(_01082_));
 sky130_fd_sc_hd__buf_4 _20716_ (.A(_04996_),
    .X(_05007_));
 sky130_fd_sc_hd__buf_4 _20717_ (.A(_03702_),
    .X(_05008_));
 sky130_fd_sc_hd__buf_4 _20718_ (.A(_04996_),
    .X(_05009_));
 sky130_fd_sc_hd__buf_12 _20719_ (.A(_12184_),
    .X(_05010_));
 sky130_fd_sc_hd__nand2_1 _20720_ (.A(_05009_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__o211a_1 _20721_ (.A1(_03222_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__mux2_1 _20722_ (.A0(_05012_),
    .A1(net3359),
    .S(_04998_),
    .X(_05013_));
 sky130_fd_sc_hd__clkbuf_1 _20723_ (.A(_05013_),
    .X(_01083_));
 sky130_fd_sc_hd__buf_12 _20724_ (.A(_12197_),
    .X(_05014_));
 sky130_fd_sc_hd__nand2_1 _20725_ (.A(_05009_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__o211a_1 _20726_ (.A1(_03228_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _20727_ (.A0(_05016_),
    .A1(net3175),
    .S(_04998_),
    .X(_05017_));
 sky130_fd_sc_hd__clkbuf_1 _20728_ (.A(_05017_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_16 _20729_ (.A(_12205_),
    .X(_05018_));
 sky130_fd_sc_hd__nand2_1 _20730_ (.A(_05009_),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__o211a_1 _20731_ (.A1(_03232_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__mux2_1 _20732_ (.A0(_05020_),
    .A1(net2441),
    .S(_04998_),
    .X(_05021_));
 sky130_fd_sc_hd__clkbuf_1 _20733_ (.A(_05021_),
    .X(_01085_));
 sky130_fd_sc_hd__buf_12 _20734_ (.A(_12213_),
    .X(_05022_));
 sky130_fd_sc_hd__nand2_1 _20735_ (.A(_05009_),
    .B(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__o211a_1 _20736_ (.A1(_03236_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__mux2_1 _20737_ (.A0(_05024_),
    .A1(net3503),
    .S(_04998_),
    .X(_05025_));
 sky130_fd_sc_hd__clkbuf_1 _20738_ (.A(_05025_),
    .X(_01086_));
 sky130_fd_sc_hd__buf_12 _20739_ (.A(_12221_),
    .X(_05026_));
 sky130_fd_sc_hd__nand2_1 _20740_ (.A(_05009_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__o211a_1 _20741_ (.A1(_03240_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__mux2_1 _20742_ (.A0(_05028_),
    .A1(net3678),
    .S(_04998_),
    .X(_05029_));
 sky130_fd_sc_hd__clkbuf_1 _20743_ (.A(_05029_),
    .X(_01087_));
 sky130_fd_sc_hd__buf_12 _20744_ (.A(_12229_),
    .X(_05030_));
 sky130_fd_sc_hd__nand2_1 _20745_ (.A(_05009_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__o211a_1 _20746_ (.A1(_03244_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__mux2_1 _20747_ (.A0(_05032_),
    .A1(net3013),
    .S(_04998_),
    .X(_05033_));
 sky130_fd_sc_hd__clkbuf_1 _20748_ (.A(_05033_),
    .X(_01088_));
 sky130_fd_sc_hd__clkbuf_16 _20749_ (.A(_12237_),
    .X(_05034_));
 sky130_fd_sc_hd__nand2_1 _20750_ (.A(_05009_),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__o211a_1 _20751_ (.A1(_03248_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_1 _20752_ (.A0(_05036_),
    .A1(net3124),
    .S(_04998_),
    .X(_05037_));
 sky130_fd_sc_hd__clkbuf_1 _20753_ (.A(_05037_),
    .X(_01089_));
 sky130_fd_sc_hd__clkbuf_16 _20754_ (.A(_12245_),
    .X(_05038_));
 sky130_fd_sc_hd__nand2_1 _20755_ (.A(_05009_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__o211a_1 _20756_ (.A1(_03252_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__mux2_1 _20757_ (.A0(_05040_),
    .A1(net2893),
    .S(_04998_),
    .X(_05041_));
 sky130_fd_sc_hd__clkbuf_1 _20758_ (.A(_05041_),
    .X(_01090_));
 sky130_fd_sc_hd__o211a_1 _20759_ (.A1(_03256_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05011_),
    .X(_05042_));
 sky130_fd_sc_hd__clkbuf_8 _20760_ (.A(_04997_),
    .X(_05043_));
 sky130_fd_sc_hd__mux2_1 _20761_ (.A0(_05042_),
    .A1(net2942),
    .S(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_1 _20762_ (.A(_05044_),
    .X(_01091_));
 sky130_fd_sc_hd__o211a_1 _20763_ (.A1(_03261_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05015_),
    .X(_05045_));
 sky130_fd_sc_hd__mux2_1 _20764_ (.A0(_05045_),
    .A1(net3402),
    .S(_05043_),
    .X(_05046_));
 sky130_fd_sc_hd__clkbuf_1 _20765_ (.A(_05046_),
    .X(_01092_));
 sky130_fd_sc_hd__o211a_1 _20766_ (.A1(_03264_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05019_),
    .X(_05047_));
 sky130_fd_sc_hd__mux2_1 _20767_ (.A0(_05047_),
    .A1(net2719),
    .S(_05043_),
    .X(_05048_));
 sky130_fd_sc_hd__clkbuf_1 _20768_ (.A(_05048_),
    .X(_01093_));
 sky130_fd_sc_hd__o211a_1 _20769_ (.A1(_03267_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05023_),
    .X(_05049_));
 sky130_fd_sc_hd__mux2_1 _20770_ (.A0(_05049_),
    .A1(net2814),
    .S(_05043_),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_1 _20771_ (.A(_05050_),
    .X(_01094_));
 sky130_fd_sc_hd__o211a_1 _20772_ (.A1(_03270_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05027_),
    .X(_05051_));
 sky130_fd_sc_hd__mux2_1 _20773_ (.A0(_05051_),
    .A1(net2512),
    .S(_05043_),
    .X(_05052_));
 sky130_fd_sc_hd__clkbuf_1 _20774_ (.A(_05052_),
    .X(_01095_));
 sky130_fd_sc_hd__o211a_1 _20775_ (.A1(_03273_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05031_),
    .X(_05053_));
 sky130_fd_sc_hd__mux2_1 _20776_ (.A0(_05053_),
    .A1(net3508),
    .S(_05043_),
    .X(_05054_));
 sky130_fd_sc_hd__clkbuf_1 _20777_ (.A(_05054_),
    .X(_01096_));
 sky130_fd_sc_hd__o211a_1 _20778_ (.A1(_03276_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05035_),
    .X(_05055_));
 sky130_fd_sc_hd__mux2_1 _20779_ (.A0(_05055_),
    .A1(net3165),
    .S(_05043_),
    .X(_05056_));
 sky130_fd_sc_hd__clkbuf_1 _20780_ (.A(_05056_),
    .X(_01097_));
 sky130_fd_sc_hd__o211a_1 _20781_ (.A1(_03279_),
    .A2(_05007_),
    .B1(_05008_),
    .C1(_05039_),
    .X(_05057_));
 sky130_fd_sc_hd__mux2_1 _20782_ (.A0(_05057_),
    .A1(net2395),
    .S(_05043_),
    .X(_05058_));
 sky130_fd_sc_hd__clkbuf_1 _20783_ (.A(_05058_),
    .X(_01098_));
 sky130_fd_sc_hd__buf_12 _20784_ (.A(_12169_),
    .X(_05059_));
 sky130_fd_sc_hd__buf_4 _20785_ (.A(_03702_),
    .X(_05060_));
 sky130_fd_sc_hd__o211a_1 _20786_ (.A1(_05059_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05011_),
    .X(_05061_));
 sky130_fd_sc_hd__mux2_1 _20787_ (.A0(_05061_),
    .A1(net3470),
    .S(_05043_),
    .X(_05062_));
 sky130_fd_sc_hd__clkbuf_1 _20788_ (.A(_05062_),
    .X(_01099_));
 sky130_fd_sc_hd__buf_12 _20789_ (.A(_12194_),
    .X(_05063_));
 sky130_fd_sc_hd__o211a_1 _20790_ (.A1(_05063_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05015_),
    .X(_05064_));
 sky130_fd_sc_hd__mux2_1 _20791_ (.A0(_05064_),
    .A1(net3033),
    .S(_05043_),
    .X(_05065_));
 sky130_fd_sc_hd__clkbuf_1 _20792_ (.A(_05065_),
    .X(_01100_));
 sky130_fd_sc_hd__clkbuf_16 _20793_ (.A(_12202_),
    .X(_05066_));
 sky130_fd_sc_hd__o211a_1 _20794_ (.A1(_05066_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05019_),
    .X(_05067_));
 sky130_fd_sc_hd__mux2_1 _20795_ (.A0(_05067_),
    .A1(net2975),
    .S(_05043_),
    .X(_05068_));
 sky130_fd_sc_hd__clkbuf_1 _20796_ (.A(_05068_),
    .X(_01101_));
 sky130_fd_sc_hd__buf_12 _20797_ (.A(_12210_),
    .X(_05069_));
 sky130_fd_sc_hd__o211a_1 _20798_ (.A1(_05069_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05023_),
    .X(_05070_));
 sky130_fd_sc_hd__mux2_1 _20799_ (.A0(_05070_),
    .A1(net2472),
    .S(_05043_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_1 _20800_ (.A(_05071_),
    .X(_01102_));
 sky130_fd_sc_hd__buf_12 _20801_ (.A(_12218_),
    .X(_05072_));
 sky130_fd_sc_hd__o211a_1 _20802_ (.A1(_05072_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05027_),
    .X(_05073_));
 sky130_fd_sc_hd__mux2_1 _20803_ (.A0(_05073_),
    .A1(net2357),
    .S(_05043_),
    .X(_05074_));
 sky130_fd_sc_hd__clkbuf_1 _20804_ (.A(_05074_),
    .X(_01103_));
 sky130_fd_sc_hd__buf_12 _20805_ (.A(_12226_),
    .X(_05075_));
 sky130_fd_sc_hd__o211a_1 _20806_ (.A1(_05075_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05031_),
    .X(_05076_));
 sky130_fd_sc_hd__mux2_1 _20807_ (.A0(_05076_),
    .A1(net2869),
    .S(_05043_),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_1 _20808_ (.A(_05077_),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_16 _20809_ (.A(_12234_),
    .X(_05078_));
 sky130_fd_sc_hd__o211a_1 _20810_ (.A1(_05078_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05035_),
    .X(_05079_));
 sky130_fd_sc_hd__mux2_1 _20811_ (.A0(_05079_),
    .A1(net3333),
    .S(_05043_),
    .X(_05080_));
 sky130_fd_sc_hd__clkbuf_1 _20812_ (.A(_05080_),
    .X(_01105_));
 sky130_fd_sc_hd__buf_12 _20813_ (.A(_12242_),
    .X(_05081_));
 sky130_fd_sc_hd__o211a_1 _20814_ (.A1(_05081_),
    .A2(_05009_),
    .B1(_05060_),
    .C1(_05039_),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _20815_ (.A0(_05082_),
    .A1(net3510),
    .S(_05043_),
    .X(_05083_));
 sky130_fd_sc_hd__clkbuf_1 _20816_ (.A(_05083_),
    .X(_01106_));
 sky130_fd_sc_hd__nand2_1 _20817_ (.A(_04995_),
    .B(_04183_),
    .Y(_05084_));
 sky130_fd_sc_hd__a21bo_1 _20818_ (.A1(_05084_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_05085_));
 sky130_fd_sc_hd__clkbuf_8 _20819_ (.A(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__mux2_1 _20820_ (.A0(_04101_),
    .A1(net3465),
    .S(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__clkbuf_1 _20821_ (.A(_05087_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _20822_ (.A0(_04109_),
    .A1(net2276),
    .S(_05086_),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _20823_ (.A(_05088_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _20824_ (.A0(_04111_),
    .A1(net2977),
    .S(_05086_),
    .X(_05089_));
 sky130_fd_sc_hd__clkbuf_1 _20825_ (.A(_05089_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _20826_ (.A0(_04113_),
    .A1(net3228),
    .S(_05086_),
    .X(_05090_));
 sky130_fd_sc_hd__clkbuf_1 _20827_ (.A(_05090_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _20828_ (.A0(_04115_),
    .A1(net2971),
    .S(_05086_),
    .X(_05091_));
 sky130_fd_sc_hd__clkbuf_1 _20829_ (.A(_05091_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _20830_ (.A0(_04117_),
    .A1(net3405),
    .S(_05086_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_1 _20831_ (.A(_05092_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _20832_ (.A0(_04119_),
    .A1(net3806),
    .S(_05086_),
    .X(_05093_));
 sky130_fd_sc_hd__clkbuf_1 _20833_ (.A(_05093_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _20834_ (.A0(_04121_),
    .A1(net3796),
    .S(_05086_),
    .X(_05094_));
 sky130_fd_sc_hd__clkbuf_1 _20835_ (.A(_05094_),
    .X(_01114_));
 sky130_fd_sc_hd__buf_12 _20836_ (.A(_02850_),
    .X(_05095_));
 sky130_fd_sc_hd__buf_4 _20837_ (.A(_05084_),
    .X(_05096_));
 sky130_fd_sc_hd__buf_4 _20838_ (.A(_05084_),
    .X(_05097_));
 sky130_fd_sc_hd__nand2_1 _20839_ (.A(_05097_),
    .B(_05010_),
    .Y(_05098_));
 sky130_fd_sc_hd__o211a_1 _20840_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__mux2_1 _20841_ (.A0(_05099_),
    .A1(net2393),
    .S(_05086_),
    .X(_05100_));
 sky130_fd_sc_hd__clkbuf_1 _20842_ (.A(_05100_),
    .X(_01115_));
 sky130_fd_sc_hd__clkbuf_16 _20843_ (.A(_02860_),
    .X(_05101_));
 sky130_fd_sc_hd__nand2_1 _20844_ (.A(_05097_),
    .B(_05014_),
    .Y(_05102_));
 sky130_fd_sc_hd__o211a_1 _20845_ (.A1(_05101_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__mux2_1 _20846_ (.A0(_05103_),
    .A1(net2557),
    .S(_05086_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_1 _20847_ (.A(_05104_),
    .X(_01116_));
 sky130_fd_sc_hd__clkbuf_16 _20848_ (.A(_02867_),
    .X(_05105_));
 sky130_fd_sc_hd__nand2_1 _20849_ (.A(_05097_),
    .B(_05018_),
    .Y(_05106_));
 sky130_fd_sc_hd__o211a_1 _20850_ (.A1(_05105_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__mux2_1 _20851_ (.A0(_05107_),
    .A1(net3520),
    .S(_05086_),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_1 _20852_ (.A(_05108_),
    .X(_01117_));
 sky130_fd_sc_hd__buf_12 _20853_ (.A(_02874_),
    .X(_05109_));
 sky130_fd_sc_hd__nand2_1 _20854_ (.A(_05097_),
    .B(_05022_),
    .Y(_05110_));
 sky130_fd_sc_hd__o211a_1 _20855_ (.A1(_05109_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__mux2_1 _20856_ (.A0(_05111_),
    .A1(net3245),
    .S(_05086_),
    .X(_05112_));
 sky130_fd_sc_hd__clkbuf_1 _20857_ (.A(_05112_),
    .X(_01118_));
 sky130_fd_sc_hd__clkbuf_16 _20858_ (.A(_02881_),
    .X(_05113_));
 sky130_fd_sc_hd__nand2_1 _20859_ (.A(_05097_),
    .B(_05026_),
    .Y(_05114_));
 sky130_fd_sc_hd__o211a_1 _20860_ (.A1(_05113_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__mux2_1 _20861_ (.A0(_05115_),
    .A1(net2856),
    .S(_05086_),
    .X(_05116_));
 sky130_fd_sc_hd__clkbuf_1 _20862_ (.A(_05116_),
    .X(_01119_));
 sky130_fd_sc_hd__clkbuf_16 _20863_ (.A(_02888_),
    .X(_05117_));
 sky130_fd_sc_hd__nand2_1 _20864_ (.A(_05097_),
    .B(_05030_),
    .Y(_05118_));
 sky130_fd_sc_hd__o211a_1 _20865_ (.A1(_05117_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__mux2_1 _20866_ (.A0(_05119_),
    .A1(net3243),
    .S(_05086_),
    .X(_05120_));
 sky130_fd_sc_hd__clkbuf_1 _20867_ (.A(_05120_),
    .X(_01120_));
 sky130_fd_sc_hd__clkbuf_16 _20868_ (.A(_02895_),
    .X(_05121_));
 sky130_fd_sc_hd__nand2_1 _20869_ (.A(_05097_),
    .B(_05034_),
    .Y(_05122_));
 sky130_fd_sc_hd__o211a_1 _20870_ (.A1(_05121_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__mux2_1 _20871_ (.A0(_05123_),
    .A1(net3058),
    .S(_05086_),
    .X(_05124_));
 sky130_fd_sc_hd__clkbuf_1 _20872_ (.A(_05124_),
    .X(_01121_));
 sky130_fd_sc_hd__clkbuf_16 _20873_ (.A(_02902_),
    .X(_05125_));
 sky130_fd_sc_hd__nand2_1 _20874_ (.A(_05097_),
    .B(_05038_),
    .Y(_05126_));
 sky130_fd_sc_hd__o211a_1 _20875_ (.A1(_05125_),
    .A2(_05096_),
    .B1(_05060_),
    .C1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _20876_ (.A0(_05127_),
    .A1(net3278),
    .S(_05086_),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _20877_ (.A(_05128_),
    .X(_01122_));
 sky130_fd_sc_hd__buf_12 _20878_ (.A(_02910_),
    .X(_05129_));
 sky130_fd_sc_hd__buf_4 _20879_ (.A(_03702_),
    .X(_05130_));
 sky130_fd_sc_hd__o211a_1 _20880_ (.A1(_05129_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05098_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_8 _20881_ (.A(_05085_),
    .X(_05132_));
 sky130_fd_sc_hd__mux2_1 _20882_ (.A0(_05131_),
    .A1(net3084),
    .S(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__clkbuf_1 _20883_ (.A(_05133_),
    .X(_01123_));
 sky130_fd_sc_hd__clkbuf_16 _20884_ (.A(_02915_),
    .X(_05134_));
 sky130_fd_sc_hd__o211a_1 _20885_ (.A1(_05134_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05102_),
    .X(_05135_));
 sky130_fd_sc_hd__mux2_1 _20886_ (.A0(_05135_),
    .A1(net3173),
    .S(_05132_),
    .X(_05136_));
 sky130_fd_sc_hd__clkbuf_1 _20887_ (.A(_05136_),
    .X(_01124_));
 sky130_fd_sc_hd__clkbuf_16 _20888_ (.A(_02920_),
    .X(_05137_));
 sky130_fd_sc_hd__o211a_1 _20889_ (.A1(_05137_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05106_),
    .X(_05138_));
 sky130_fd_sc_hd__mux2_1 _20890_ (.A0(_05138_),
    .A1(net3502),
    .S(_05132_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_1 _20891_ (.A(_05139_),
    .X(_01125_));
 sky130_fd_sc_hd__buf_12 _20892_ (.A(_02926_),
    .X(_05140_));
 sky130_fd_sc_hd__o211a_1 _20893_ (.A1(_05140_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05110_),
    .X(_05141_));
 sky130_fd_sc_hd__mux2_1 _20894_ (.A0(_05141_),
    .A1(net3318),
    .S(_05132_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_1 _20895_ (.A(_05142_),
    .X(_01126_));
 sky130_fd_sc_hd__clkbuf_16 _20896_ (.A(_02931_),
    .X(_05143_));
 sky130_fd_sc_hd__o211a_1 _20897_ (.A1(_05143_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05114_),
    .X(_05144_));
 sky130_fd_sc_hd__mux2_1 _20898_ (.A0(_05144_),
    .A1(net2747),
    .S(_05132_),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_1 _20899_ (.A(_05145_),
    .X(_01127_));
 sky130_fd_sc_hd__buf_12 _20900_ (.A(_02936_),
    .X(_05146_));
 sky130_fd_sc_hd__o211a_1 _20901_ (.A1(_05146_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05118_),
    .X(_05147_));
 sky130_fd_sc_hd__mux2_1 _20902_ (.A0(_05147_),
    .A1(net3148),
    .S(_05132_),
    .X(_05148_));
 sky130_fd_sc_hd__clkbuf_1 _20903_ (.A(_05148_),
    .X(_01128_));
 sky130_fd_sc_hd__clkbuf_16 _20904_ (.A(_02941_),
    .X(_05149_));
 sky130_fd_sc_hd__o211a_1 _20905_ (.A1(_05149_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05122_),
    .X(_05150_));
 sky130_fd_sc_hd__mux2_1 _20906_ (.A0(_05150_),
    .A1(net3562),
    .S(_05132_),
    .X(_05151_));
 sky130_fd_sc_hd__clkbuf_1 _20907_ (.A(_05151_),
    .X(_01129_));
 sky130_fd_sc_hd__buf_8 _20908_ (.A(_02946_),
    .X(_05152_));
 sky130_fd_sc_hd__o211a_1 _20909_ (.A1(_05152_),
    .A2(_05096_),
    .B1(_05130_),
    .C1(_05126_),
    .X(_05153_));
 sky130_fd_sc_hd__mux2_1 _20910_ (.A0(_05153_),
    .A1(net3346),
    .S(_05132_),
    .X(_05154_));
 sky130_fd_sc_hd__clkbuf_1 _20911_ (.A(_05154_),
    .X(_01130_));
 sky130_fd_sc_hd__o211a_1 _20912_ (.A1(_05059_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05098_),
    .X(_05155_));
 sky130_fd_sc_hd__mux2_1 _20913_ (.A0(_05155_),
    .A1(net3217),
    .S(_05132_),
    .X(_05156_));
 sky130_fd_sc_hd__clkbuf_1 _20914_ (.A(_05156_),
    .X(_01131_));
 sky130_fd_sc_hd__o211a_1 _20915_ (.A1(_05063_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05102_),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_1 _20916_ (.A0(_05157_),
    .A1(net2759),
    .S(_05132_),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_1 _20917_ (.A(_05158_),
    .X(_01132_));
 sky130_fd_sc_hd__o211a_1 _20918_ (.A1(_05066_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05106_),
    .X(_05159_));
 sky130_fd_sc_hd__mux2_1 _20919_ (.A0(_05159_),
    .A1(net3528),
    .S(_05132_),
    .X(_05160_));
 sky130_fd_sc_hd__clkbuf_1 _20920_ (.A(_05160_),
    .X(_01133_));
 sky130_fd_sc_hd__o211a_1 _20921_ (.A1(_05069_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05110_),
    .X(_05161_));
 sky130_fd_sc_hd__mux2_1 _20922_ (.A0(_05161_),
    .A1(net2379),
    .S(_05132_),
    .X(_05162_));
 sky130_fd_sc_hd__clkbuf_1 _20923_ (.A(_05162_),
    .X(_01134_));
 sky130_fd_sc_hd__o211a_1 _20924_ (.A1(_05072_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05114_),
    .X(_05163_));
 sky130_fd_sc_hd__mux2_1 _20925_ (.A0(_05163_),
    .A1(net3233),
    .S(_05132_),
    .X(_05164_));
 sky130_fd_sc_hd__clkbuf_1 _20926_ (.A(_05164_),
    .X(_01135_));
 sky130_fd_sc_hd__o211a_1 _20927_ (.A1(_05075_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05118_),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_1 _20928_ (.A0(_05165_),
    .A1(net2790),
    .S(_05132_),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _20929_ (.A(_05166_),
    .X(_01136_));
 sky130_fd_sc_hd__o211a_1 _20930_ (.A1(_05078_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05122_),
    .X(_05167_));
 sky130_fd_sc_hd__mux2_1 _20931_ (.A0(_05167_),
    .A1(net3206),
    .S(_05132_),
    .X(_05168_));
 sky130_fd_sc_hd__clkbuf_1 _20932_ (.A(_05168_),
    .X(_01137_));
 sky130_fd_sc_hd__o211a_1 _20933_ (.A1(_05081_),
    .A2(_05097_),
    .B1(_05130_),
    .C1(_05126_),
    .X(_05169_));
 sky130_fd_sc_hd__mux2_1 _20934_ (.A0(_05169_),
    .A1(net3695),
    .S(_05132_),
    .X(_05170_));
 sky130_fd_sc_hd__clkbuf_1 _20935_ (.A(_05170_),
    .X(_01138_));
 sky130_fd_sc_hd__nand2_1 _20936_ (.A(_04995_),
    .B(_04257_),
    .Y(_05171_));
 sky130_fd_sc_hd__a21bo_1 _20937_ (.A1(_05171_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_05172_));
 sky130_fd_sc_hd__buf_6 _20938_ (.A(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__mux2_1 _20939_ (.A0(_04101_),
    .A1(net3549),
    .S(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__clkbuf_1 _20940_ (.A(_05174_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _20941_ (.A0(_04109_),
    .A1(net2846),
    .S(_05173_),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_1 _20942_ (.A(_05175_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _20943_ (.A0(_04111_),
    .A1(net2401),
    .S(_05173_),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_1 _20944_ (.A(_05176_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _20945_ (.A0(_04113_),
    .A1(net2940),
    .S(_05173_),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_1 _20946_ (.A(_05177_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _20947_ (.A0(_04115_),
    .A1(net3430),
    .S(_05173_),
    .X(_05178_));
 sky130_fd_sc_hd__clkbuf_1 _20948_ (.A(_05178_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _20949_ (.A0(_04117_),
    .A1(net3227),
    .S(_05173_),
    .X(_05179_));
 sky130_fd_sc_hd__clkbuf_1 _20950_ (.A(_05179_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _20951_ (.A0(_04119_),
    .A1(net3839),
    .S(_05173_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_1 _20952_ (.A(_05180_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _20953_ (.A0(_04121_),
    .A1(net3729),
    .S(_05173_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _20954_ (.A(_05181_),
    .X(_01146_));
 sky130_fd_sc_hd__buf_4 _20955_ (.A(_05171_),
    .X(_05182_));
 sky130_fd_sc_hd__buf_8 _20956_ (.A(_09125_),
    .X(_05183_));
 sky130_fd_sc_hd__buf_4 _20957_ (.A(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__buf_4 _20958_ (.A(_05171_),
    .X(_05185_));
 sky130_fd_sc_hd__nand2_1 _20959_ (.A(_05185_),
    .B(_05010_),
    .Y(_05186_));
 sky130_fd_sc_hd__o211a_1 _20960_ (.A1(_05095_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_1 _20961_ (.A0(_05187_),
    .A1(net3120),
    .S(_05173_),
    .X(_05188_));
 sky130_fd_sc_hd__clkbuf_1 _20962_ (.A(_05188_),
    .X(_01147_));
 sky130_fd_sc_hd__nand2_1 _20963_ (.A(_05185_),
    .B(_05014_),
    .Y(_05189_));
 sky130_fd_sc_hd__o211a_1 _20964_ (.A1(_05101_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__mux2_1 _20965_ (.A0(_05190_),
    .A1(net2118),
    .S(_05173_),
    .X(_05191_));
 sky130_fd_sc_hd__clkbuf_1 _20966_ (.A(_05191_),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _20967_ (.A(_05185_),
    .B(_05018_),
    .Y(_05192_));
 sky130_fd_sc_hd__o211a_1 _20968_ (.A1(_05105_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__mux2_1 _20969_ (.A0(_05193_),
    .A1(net3464),
    .S(_05173_),
    .X(_05194_));
 sky130_fd_sc_hd__clkbuf_1 _20970_ (.A(_05194_),
    .X(_01149_));
 sky130_fd_sc_hd__nand2_1 _20971_ (.A(_05185_),
    .B(_05022_),
    .Y(_05195_));
 sky130_fd_sc_hd__o211a_1 _20972_ (.A1(_05109_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _20973_ (.A0(_05196_),
    .A1(net2838),
    .S(_05173_),
    .X(_05197_));
 sky130_fd_sc_hd__clkbuf_1 _20974_ (.A(_05197_),
    .X(_01150_));
 sky130_fd_sc_hd__nand2_1 _20975_ (.A(_05185_),
    .B(_05026_),
    .Y(_05198_));
 sky130_fd_sc_hd__o211a_1 _20976_ (.A1(_05113_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_1 _20977_ (.A0(_05199_),
    .A1(net2124),
    .S(_05173_),
    .X(_05200_));
 sky130_fd_sc_hd__clkbuf_1 _20978_ (.A(_05200_),
    .X(_01151_));
 sky130_fd_sc_hd__nand2_1 _20979_ (.A(_05185_),
    .B(_05030_),
    .Y(_05201_));
 sky130_fd_sc_hd__o211a_1 _20980_ (.A1(_05117_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__mux2_1 _20981_ (.A0(_05202_),
    .A1(net2184),
    .S(_05173_),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_1 _20982_ (.A(_05203_),
    .X(_01152_));
 sky130_fd_sc_hd__nand2_1 _20983_ (.A(_05185_),
    .B(_05034_),
    .Y(_05204_));
 sky130_fd_sc_hd__o211a_1 _20984_ (.A1(_05121_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__mux2_1 _20985_ (.A0(_05205_),
    .A1(net3053),
    .S(_05173_),
    .X(_05206_));
 sky130_fd_sc_hd__clkbuf_1 _20986_ (.A(_05206_),
    .X(_01153_));
 sky130_fd_sc_hd__nand2_1 _20987_ (.A(_05185_),
    .B(_05038_),
    .Y(_05207_));
 sky130_fd_sc_hd__o211a_1 _20988_ (.A1(_05125_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__mux2_1 _20989_ (.A0(_05208_),
    .A1(net3032),
    .S(_05173_),
    .X(_05209_));
 sky130_fd_sc_hd__clkbuf_1 _20990_ (.A(_05209_),
    .X(_01154_));
 sky130_fd_sc_hd__o211a_1 _20991_ (.A1(_05129_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05186_),
    .X(_05210_));
 sky130_fd_sc_hd__clkbuf_8 _20992_ (.A(_05172_),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_1 _20993_ (.A0(_05210_),
    .A1(net3162),
    .S(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_1 _20994_ (.A(_05212_),
    .X(_01155_));
 sky130_fd_sc_hd__o211a_1 _20995_ (.A1(_05134_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05189_),
    .X(_05213_));
 sky130_fd_sc_hd__mux2_1 _20996_ (.A0(_05213_),
    .A1(net3209),
    .S(_05211_),
    .X(_05214_));
 sky130_fd_sc_hd__clkbuf_1 _20997_ (.A(_05214_),
    .X(_01156_));
 sky130_fd_sc_hd__o211a_1 _20998_ (.A1(_05137_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05192_),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _20999_ (.A0(_05215_),
    .A1(net2886),
    .S(_05211_),
    .X(_05216_));
 sky130_fd_sc_hd__clkbuf_1 _21000_ (.A(_05216_),
    .X(_01157_));
 sky130_fd_sc_hd__o211a_1 _21001_ (.A1(_05140_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05195_),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_1 _21002_ (.A0(_05217_),
    .A1(net3596),
    .S(_05211_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_1 _21003_ (.A(_05218_),
    .X(_01158_));
 sky130_fd_sc_hd__o211a_1 _21004_ (.A1(_05143_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05198_),
    .X(_05219_));
 sky130_fd_sc_hd__mux2_1 _21005_ (.A0(_05219_),
    .A1(net3450),
    .S(_05211_),
    .X(_05220_));
 sky130_fd_sc_hd__clkbuf_1 _21006_ (.A(_05220_),
    .X(_01159_));
 sky130_fd_sc_hd__o211a_1 _21007_ (.A1(_05146_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05201_),
    .X(_05221_));
 sky130_fd_sc_hd__mux2_1 _21008_ (.A0(_05221_),
    .A1(net3052),
    .S(_05211_),
    .X(_05222_));
 sky130_fd_sc_hd__clkbuf_1 _21009_ (.A(_05222_),
    .X(_01160_));
 sky130_fd_sc_hd__o211a_1 _21010_ (.A1(_05149_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05204_),
    .X(_05223_));
 sky130_fd_sc_hd__mux2_1 _21011_ (.A0(_05223_),
    .A1(net3517),
    .S(_05211_),
    .X(_05224_));
 sky130_fd_sc_hd__clkbuf_1 _21012_ (.A(_05224_),
    .X(_01161_));
 sky130_fd_sc_hd__o211a_1 _21013_ (.A1(_05152_),
    .A2(_05182_),
    .B1(_05184_),
    .C1(_05207_),
    .X(_05225_));
 sky130_fd_sc_hd__mux2_1 _21014_ (.A0(_05225_),
    .A1(net3543),
    .S(_05211_),
    .X(_05226_));
 sky130_fd_sc_hd__clkbuf_1 _21015_ (.A(_05226_),
    .X(_01162_));
 sky130_fd_sc_hd__buf_4 _21016_ (.A(_05183_),
    .X(_05227_));
 sky130_fd_sc_hd__o211a_1 _21017_ (.A1(_05059_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05186_),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _21018_ (.A0(_05228_),
    .A1(net2986),
    .S(_05211_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_1 _21019_ (.A(_05229_),
    .X(_01163_));
 sky130_fd_sc_hd__o211a_1 _21020_ (.A1(_05063_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05189_),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _21021_ (.A0(_05230_),
    .A1(net2934),
    .S(_05211_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _21022_ (.A(_05231_),
    .X(_01164_));
 sky130_fd_sc_hd__o211a_1 _21023_ (.A1(_05066_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05192_),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _21024_ (.A0(_05232_),
    .A1(net2717),
    .S(_05211_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _21025_ (.A(_05233_),
    .X(_01165_));
 sky130_fd_sc_hd__o211a_1 _21026_ (.A1(_05069_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05195_),
    .X(_05234_));
 sky130_fd_sc_hd__mux2_1 _21027_ (.A0(_05234_),
    .A1(net2962),
    .S(_05211_),
    .X(_05235_));
 sky130_fd_sc_hd__clkbuf_1 _21028_ (.A(_05235_),
    .X(_01166_));
 sky130_fd_sc_hd__o211a_1 _21029_ (.A1(_05072_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05198_),
    .X(_05236_));
 sky130_fd_sc_hd__mux2_1 _21030_ (.A0(_05236_),
    .A1(net2281),
    .S(_05211_),
    .X(_05237_));
 sky130_fd_sc_hd__clkbuf_1 _21031_ (.A(_05237_),
    .X(_01167_));
 sky130_fd_sc_hd__o211a_1 _21032_ (.A1(_05075_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05201_),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_1 _21033_ (.A0(_05238_),
    .A1(net3019),
    .S(_05211_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_1 _21034_ (.A(_05239_),
    .X(_01168_));
 sky130_fd_sc_hd__o211a_1 _21035_ (.A1(_05078_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05204_),
    .X(_05240_));
 sky130_fd_sc_hd__mux2_1 _21036_ (.A0(_05240_),
    .A1(net3224),
    .S(_05211_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _21037_ (.A(_05241_),
    .X(_01169_));
 sky130_fd_sc_hd__o211a_1 _21038_ (.A1(_05081_),
    .A2(_05185_),
    .B1(_05227_),
    .C1(_05207_),
    .X(_05242_));
 sky130_fd_sc_hd__mux2_1 _21039_ (.A0(_05242_),
    .A1(net2207),
    .S(_05211_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_1 _21040_ (.A(_05243_),
    .X(_01170_));
 sky130_fd_sc_hd__nand2_1 _21041_ (.A(_04995_),
    .B(_04333_),
    .Y(_05244_));
 sky130_fd_sc_hd__inv_2 _21042_ (.A(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__o21ai_4 _21043_ (.A1(_04332_),
    .A2(_05245_),
    .B1(_04776_),
    .Y(_05246_));
 sky130_fd_sc_hd__mux2_1 _21044_ (.A0(_04101_),
    .A1(net3045),
    .S(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__clkbuf_1 _21045_ (.A(_05247_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _21046_ (.A0(_04109_),
    .A1(net2519),
    .S(_05246_),
    .X(_05248_));
 sky130_fd_sc_hd__clkbuf_1 _21047_ (.A(_05248_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _21048_ (.A0(_04111_),
    .A1(net2780),
    .S(_05246_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _21049_ (.A(_05249_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _21050_ (.A0(_04113_),
    .A1(net2899),
    .S(_05246_),
    .X(_05250_));
 sky130_fd_sc_hd__clkbuf_1 _21051_ (.A(_05250_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _21052_ (.A0(_04115_),
    .A1(net3030),
    .S(_05246_),
    .X(_05251_));
 sky130_fd_sc_hd__clkbuf_1 _21053_ (.A(_05251_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _21054_ (.A0(_04117_),
    .A1(net2807),
    .S(_05246_),
    .X(_05252_));
 sky130_fd_sc_hd__clkbuf_1 _21055_ (.A(_05252_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _21056_ (.A0(_04119_),
    .A1(net2684),
    .S(_05246_),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_1 _21057_ (.A(_05253_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _21058_ (.A0(_04121_),
    .A1(net3499),
    .S(_05246_),
    .X(_05254_));
 sky130_fd_sc_hd__clkbuf_1 _21059_ (.A(_05254_),
    .X(_01178_));
 sky130_fd_sc_hd__buf_4 _21060_ (.A(_05246_),
    .X(_05255_));
 sky130_fd_sc_hd__buf_4 _21061_ (.A(_05245_),
    .X(_05256_));
 sky130_fd_sc_hd__buf_4 _21062_ (.A(_05245_),
    .X(_05257_));
 sky130_fd_sc_hd__nor2_1 _21063_ (.A(_02854_),
    .B(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__a211o_1 _21064_ (.A1(_02852_),
    .A2(_05256_),
    .B1(_04966_),
    .C1(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__buf_4 _21065_ (.A(_05246_),
    .X(_05260_));
 sky130_fd_sc_hd__nand2_1 _21066_ (.A(_05260_),
    .B(net1294),
    .Y(_05261_));
 sky130_fd_sc_hd__o21ai_1 _21067_ (.A1(_05255_),
    .A2(_05259_),
    .B1(net1295),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _21068_ (.A(_02863_),
    .B(_05257_),
    .Y(_05262_));
 sky130_fd_sc_hd__a211o_1 _21069_ (.A1(_02862_),
    .A2(_05256_),
    .B1(_04966_),
    .C1(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__nand2_1 _21070_ (.A(_05260_),
    .B(net1164),
    .Y(_05264_));
 sky130_fd_sc_hd__o21ai_1 _21071_ (.A1(_05255_),
    .A2(_05263_),
    .B1(net1165),
    .Y(_01180_));
 sky130_fd_sc_hd__buf_4 _21072_ (.A(_04598_),
    .X(_05265_));
 sky130_fd_sc_hd__nor2_1 _21073_ (.A(_02870_),
    .B(_05257_),
    .Y(_05266_));
 sky130_fd_sc_hd__a211o_1 _21074_ (.A1(_02869_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__nand2_1 _21075_ (.A(_05260_),
    .B(net1162),
    .Y(_05268_));
 sky130_fd_sc_hd__o21ai_1 _21076_ (.A1(_05255_),
    .A2(_05267_),
    .B1(net1163),
    .Y(_01181_));
 sky130_fd_sc_hd__nor2_1 _21077_ (.A(_02877_),
    .B(_05257_),
    .Y(_05269_));
 sky130_fd_sc_hd__a211o_1 _21078_ (.A1(_02876_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__nand2_1 _21079_ (.A(_05260_),
    .B(net528),
    .Y(_05271_));
 sky130_fd_sc_hd__o21ai_1 _21080_ (.A1(_05255_),
    .A2(_05270_),
    .B1(net529),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _21081_ (.A(_02884_),
    .B(_05257_),
    .Y(_05272_));
 sky130_fd_sc_hd__a211o_1 _21082_ (.A1(_02883_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__nand2_1 _21083_ (.A(_05260_),
    .B(net694),
    .Y(_05274_));
 sky130_fd_sc_hd__o21ai_1 _21084_ (.A1(_05255_),
    .A2(_05273_),
    .B1(net695),
    .Y(_01183_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(_02891_),
    .B(_05257_),
    .Y(_05275_));
 sky130_fd_sc_hd__a211o_1 _21086_ (.A1(_02890_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__nand2_1 _21087_ (.A(_05260_),
    .B(net578),
    .Y(_05277_));
 sky130_fd_sc_hd__o21ai_1 _21088_ (.A1(_05255_),
    .A2(_05276_),
    .B1(net579),
    .Y(_01184_));
 sky130_fd_sc_hd__nor2_1 _21089_ (.A(_02898_),
    .B(_05257_),
    .Y(_05278_));
 sky130_fd_sc_hd__a211o_1 _21090_ (.A1(_02897_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__nand2_1 _21091_ (.A(_05260_),
    .B(net772),
    .Y(_05280_));
 sky130_fd_sc_hd__o21ai_1 _21092_ (.A1(_05255_),
    .A2(_05279_),
    .B1(net773),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _21093_ (.A(_02905_),
    .B(_05257_),
    .Y(_05281_));
 sky130_fd_sc_hd__a211o_1 _21094_ (.A1(_02904_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__nand2_1 _21095_ (.A(_05260_),
    .B(net1520),
    .Y(_05283_));
 sky130_fd_sc_hd__o21ai_1 _21096_ (.A1(_05255_),
    .A2(_05282_),
    .B1(net1521),
    .Y(_01186_));
 sky130_fd_sc_hd__buf_4 _21097_ (.A(_05246_),
    .X(_05284_));
 sky130_fd_sc_hd__a211o_1 _21098_ (.A1(_02912_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05258_),
    .X(_05285_));
 sky130_fd_sc_hd__nand2_1 _21099_ (.A(_05260_),
    .B(net1228),
    .Y(_05286_));
 sky130_fd_sc_hd__o21ai_1 _21100_ (.A1(_05284_),
    .A2(_05285_),
    .B1(net1229),
    .Y(_01187_));
 sky130_fd_sc_hd__a211o_1 _21101_ (.A1(_02917_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05262_),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _21102_ (.A(_05260_),
    .B(net1674),
    .Y(_05288_));
 sky130_fd_sc_hd__o21ai_1 _21103_ (.A1(_05284_),
    .A2(_05287_),
    .B1(net1675),
    .Y(_01188_));
 sky130_fd_sc_hd__a211o_1 _21104_ (.A1(_02922_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05266_),
    .X(_05289_));
 sky130_fd_sc_hd__nand2_1 _21105_ (.A(_05260_),
    .B(net1110),
    .Y(_05290_));
 sky130_fd_sc_hd__o21ai_1 _21106_ (.A1(_05284_),
    .A2(_05289_),
    .B1(net1111),
    .Y(_01189_));
 sky130_fd_sc_hd__a211o_1 _21107_ (.A1(_02928_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05269_),
    .X(_05291_));
 sky130_fd_sc_hd__nand2_1 _21108_ (.A(_05260_),
    .B(net930),
    .Y(_05292_));
 sky130_fd_sc_hd__o21ai_1 _21109_ (.A1(_05284_),
    .A2(_05291_),
    .B1(net931),
    .Y(_01190_));
 sky130_fd_sc_hd__a211o_1 _21110_ (.A1(_02933_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05272_),
    .X(_05293_));
 sky130_fd_sc_hd__nand2_1 _21111_ (.A(_05260_),
    .B(net1062),
    .Y(_05294_));
 sky130_fd_sc_hd__o21ai_1 _21112_ (.A1(_05284_),
    .A2(_05293_),
    .B1(net1063),
    .Y(_01191_));
 sky130_fd_sc_hd__a211o_1 _21113_ (.A1(_02938_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05275_),
    .X(_05295_));
 sky130_fd_sc_hd__nand2_1 _21114_ (.A(_05260_),
    .B(net1006),
    .Y(_05296_));
 sky130_fd_sc_hd__o21ai_1 _21115_ (.A1(_05284_),
    .A2(_05295_),
    .B1(net1007),
    .Y(_01192_));
 sky130_fd_sc_hd__a211o_1 _21116_ (.A1(_02943_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05278_),
    .X(_05297_));
 sky130_fd_sc_hd__nand2_1 _21117_ (.A(_05260_),
    .B(net1584),
    .Y(_05298_));
 sky130_fd_sc_hd__o21ai_1 _21118_ (.A1(_05284_),
    .A2(_05297_),
    .B1(net1585),
    .Y(_01193_));
 sky130_fd_sc_hd__a211o_1 _21119_ (.A1(_02948_),
    .A2(_05256_),
    .B1(_05265_),
    .C1(_05281_),
    .X(_05299_));
 sky130_fd_sc_hd__nand2_1 _21120_ (.A(_05260_),
    .B(net1154),
    .Y(_05300_));
 sky130_fd_sc_hd__o21ai_1 _21121_ (.A1(_05284_),
    .A2(_05299_),
    .B1(net1155),
    .Y(_01194_));
 sky130_fd_sc_hd__a211o_1 _21122_ (.A1(_02952_),
    .A2(_05257_),
    .B1(_05265_),
    .C1(_05258_),
    .X(_05301_));
 sky130_fd_sc_hd__nand2_1 _21123_ (.A(_05255_),
    .B(net1710),
    .Y(_05302_));
 sky130_fd_sc_hd__o21ai_1 _21124_ (.A1(_05284_),
    .A2(_05301_),
    .B1(net1711),
    .Y(_01195_));
 sky130_fd_sc_hd__a211o_1 _21125_ (.A1(_02956_),
    .A2(_05257_),
    .B1(_05265_),
    .C1(_05262_),
    .X(_05303_));
 sky130_fd_sc_hd__nand2_1 _21126_ (.A(_05255_),
    .B(net1700),
    .Y(_05304_));
 sky130_fd_sc_hd__o21ai_1 _21127_ (.A1(_05284_),
    .A2(_05303_),
    .B1(net1701),
    .Y(_01196_));
 sky130_fd_sc_hd__buf_4 _21128_ (.A(_04598_),
    .X(_05305_));
 sky130_fd_sc_hd__a211o_1 _21129_ (.A1(_02960_),
    .A2(_05257_),
    .B1(_05305_),
    .C1(_05266_),
    .X(_05306_));
 sky130_fd_sc_hd__nand2_1 _21130_ (.A(_05255_),
    .B(net1234),
    .Y(_05307_));
 sky130_fd_sc_hd__o21ai_1 _21131_ (.A1(_05284_),
    .A2(_05306_),
    .B1(net1235),
    .Y(_01197_));
 sky130_fd_sc_hd__a211o_1 _21132_ (.A1(_02964_),
    .A2(_05257_),
    .B1(_05305_),
    .C1(_05269_),
    .X(_05308_));
 sky130_fd_sc_hd__nand2_1 _21133_ (.A(_05255_),
    .B(net1178),
    .Y(_05309_));
 sky130_fd_sc_hd__o21ai_1 _21134_ (.A1(_05284_),
    .A2(_05308_),
    .B1(net1179),
    .Y(_01198_));
 sky130_fd_sc_hd__a211o_1 _21135_ (.A1(_02968_),
    .A2(_05257_),
    .B1(_05305_),
    .C1(_05272_),
    .X(_05310_));
 sky130_fd_sc_hd__nand2_1 _21136_ (.A(_05255_),
    .B(net1338),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_1 _21137_ (.A1(_05284_),
    .A2(_05310_),
    .B1(net1339),
    .Y(_01199_));
 sky130_fd_sc_hd__a211o_1 _21138_ (.A1(_02972_),
    .A2(_05257_),
    .B1(_05305_),
    .C1(_05275_),
    .X(_05312_));
 sky130_fd_sc_hd__nand2_1 _21139_ (.A(_05255_),
    .B(net1438),
    .Y(_05313_));
 sky130_fd_sc_hd__o21ai_1 _21140_ (.A1(_05284_),
    .A2(_05312_),
    .B1(net1439),
    .Y(_01200_));
 sky130_fd_sc_hd__a211o_1 _21141_ (.A1(_02976_),
    .A2(_05257_),
    .B1(_05305_),
    .C1(_05278_),
    .X(_05314_));
 sky130_fd_sc_hd__nand2_1 _21142_ (.A(_05255_),
    .B(net1140),
    .Y(_05315_));
 sky130_fd_sc_hd__o21ai_1 _21143_ (.A1(_05284_),
    .A2(_05314_),
    .B1(net1141),
    .Y(_01201_));
 sky130_fd_sc_hd__a211o_1 _21144_ (.A1(_02980_),
    .A2(_05257_),
    .B1(_05305_),
    .C1(_05281_),
    .X(_05316_));
 sky130_fd_sc_hd__nand2_1 _21145_ (.A(_05255_),
    .B(net816),
    .Y(_05317_));
 sky130_fd_sc_hd__o21ai_1 _21146_ (.A1(_05284_),
    .A2(_05316_),
    .B1(net817),
    .Y(_01202_));
 sky130_fd_sc_hd__buf_8 _21147_ (.A(_02809_),
    .X(_05318_));
 sky130_fd_sc_hd__and3_4 _21148_ (.A(_02813_),
    .B(\line_cache_idx[7] ),
    .C(_12303_),
    .X(_05319_));
 sky130_fd_sc_hd__nand2_1 _21149_ (.A(_05319_),
    .B(_04104_),
    .Y(_05320_));
 sky130_fd_sc_hd__a21bo_1 _21150_ (.A1(_05320_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_8 _21151_ (.A(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__mux2_1 _21152_ (.A0(_05318_),
    .A1(net2044),
    .S(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_1 _21153_ (.A(_05323_),
    .X(_01203_));
 sky130_fd_sc_hd__buf_12 _21154_ (.A(_02822_),
    .X(_05324_));
 sky130_fd_sc_hd__mux2_1 _21155_ (.A0(_05324_),
    .A1(net2520),
    .S(_05322_),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _21156_ (.A(_05325_),
    .X(_01204_));
 sky130_fd_sc_hd__clkbuf_16 _21157_ (.A(_02826_),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_1 _21158_ (.A0(_05326_),
    .A1(net2093),
    .S(_05322_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _21159_ (.A(_05327_),
    .X(_01205_));
 sky130_fd_sc_hd__buf_8 _21160_ (.A(_02830_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_1 _21161_ (.A0(_05328_),
    .A1(net3067),
    .S(_05322_),
    .X(_05329_));
 sky130_fd_sc_hd__clkbuf_1 _21162_ (.A(_05329_),
    .X(_01206_));
 sky130_fd_sc_hd__clkbuf_16 _21163_ (.A(_02834_),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_1 _21164_ (.A0(_05330_),
    .A1(net3070),
    .S(_05322_),
    .X(_05331_));
 sky130_fd_sc_hd__clkbuf_1 _21165_ (.A(_05331_),
    .X(_01207_));
 sky130_fd_sc_hd__buf_8 _21166_ (.A(_02838_),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_1 _21167_ (.A0(_05332_),
    .A1(net3573),
    .S(_05322_),
    .X(_05333_));
 sky130_fd_sc_hd__clkbuf_1 _21168_ (.A(_05333_),
    .X(_01208_));
 sky130_fd_sc_hd__buf_8 _21169_ (.A(_02842_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _21170_ (.A0(_05334_),
    .A1(net2575),
    .S(_05322_),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _21171_ (.A(_05335_),
    .X(_01209_));
 sky130_fd_sc_hd__buf_8 _21172_ (.A(_02846_),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _21173_ (.A0(_05336_),
    .A1(net2069),
    .S(_05322_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _21174_ (.A(_05337_),
    .X(_01210_));
 sky130_fd_sc_hd__buf_4 _21175_ (.A(_05320_),
    .X(_05338_));
 sky130_fd_sc_hd__buf_4 _21176_ (.A(_05320_),
    .X(_05339_));
 sky130_fd_sc_hd__nand2_1 _21177_ (.A(_05339_),
    .B(_05010_),
    .Y(_05340_));
 sky130_fd_sc_hd__o211a_1 _21178_ (.A1(_05095_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__mux2_1 _21179_ (.A0(_05341_),
    .A1(net2833),
    .S(_05322_),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_1 _21180_ (.A(_05342_),
    .X(_01211_));
 sky130_fd_sc_hd__nand2_1 _21181_ (.A(_05339_),
    .B(_05014_),
    .Y(_05343_));
 sky130_fd_sc_hd__o211a_1 _21182_ (.A1(_05101_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_1 _21183_ (.A0(_05344_),
    .A1(net2896),
    .S(_05322_),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _21184_ (.A(_05345_),
    .X(_01212_));
 sky130_fd_sc_hd__nand2_1 _21185_ (.A(_05339_),
    .B(_05018_),
    .Y(_05346_));
 sky130_fd_sc_hd__o211a_1 _21186_ (.A1(_05105_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__mux2_1 _21187_ (.A0(_05347_),
    .A1(net3121),
    .S(_05322_),
    .X(_05348_));
 sky130_fd_sc_hd__clkbuf_1 _21188_ (.A(_05348_),
    .X(_01213_));
 sky130_fd_sc_hd__nand2_1 _21189_ (.A(_05339_),
    .B(_05022_),
    .Y(_05349_));
 sky130_fd_sc_hd__o211a_1 _21190_ (.A1(_05109_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__mux2_1 _21191_ (.A0(_05350_),
    .A1(net3383),
    .S(_05322_),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _21192_ (.A(_05351_),
    .X(_01214_));
 sky130_fd_sc_hd__nand2_1 _21193_ (.A(_05339_),
    .B(_05026_),
    .Y(_05352_));
 sky130_fd_sc_hd__o211a_1 _21194_ (.A1(_05113_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__mux2_1 _21195_ (.A0(_05353_),
    .A1(net3330),
    .S(_05322_),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_1 _21196_ (.A(_05354_),
    .X(_01215_));
 sky130_fd_sc_hd__nand2_1 _21197_ (.A(_05339_),
    .B(_05030_),
    .Y(_05355_));
 sky130_fd_sc_hd__o211a_1 _21198_ (.A1(_05117_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__mux2_1 _21199_ (.A0(_05356_),
    .A1(net2589),
    .S(_05322_),
    .X(_05357_));
 sky130_fd_sc_hd__clkbuf_1 _21200_ (.A(_05357_),
    .X(_01216_));
 sky130_fd_sc_hd__nand2_1 _21201_ (.A(_05339_),
    .B(_05034_),
    .Y(_05358_));
 sky130_fd_sc_hd__o211a_1 _21202_ (.A1(_05121_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__mux2_1 _21203_ (.A0(_05359_),
    .A1(net2961),
    .S(_05322_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _21204_ (.A(_05360_),
    .X(_01217_));
 sky130_fd_sc_hd__nand2_1 _21205_ (.A(_05339_),
    .B(_05038_),
    .Y(_05361_));
 sky130_fd_sc_hd__o211a_1 _21206_ (.A1(_05125_),
    .A2(_05338_),
    .B1(_05227_),
    .C1(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__mux2_1 _21207_ (.A0(_05362_),
    .A1(net2658),
    .S(_05322_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _21208_ (.A(_05363_),
    .X(_01218_));
 sky130_fd_sc_hd__buf_4 _21209_ (.A(_05183_),
    .X(_05364_));
 sky130_fd_sc_hd__o211a_1 _21210_ (.A1(_05129_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05340_),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_8 _21211_ (.A(_05321_),
    .X(_05366_));
 sky130_fd_sc_hd__mux2_1 _21212_ (.A0(_05365_),
    .A1(net3213),
    .S(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _21213_ (.A(_05367_),
    .X(_01219_));
 sky130_fd_sc_hd__o211a_1 _21214_ (.A1(_05134_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05343_),
    .X(_05368_));
 sky130_fd_sc_hd__mux2_1 _21215_ (.A0(_05368_),
    .A1(net3117),
    .S(_05366_),
    .X(_05369_));
 sky130_fd_sc_hd__clkbuf_1 _21216_ (.A(_05369_),
    .X(_01220_));
 sky130_fd_sc_hd__o211a_1 _21217_ (.A1(_05137_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05346_),
    .X(_05370_));
 sky130_fd_sc_hd__mux2_1 _21218_ (.A0(_05370_),
    .A1(net3522),
    .S(_05366_),
    .X(_05371_));
 sky130_fd_sc_hd__clkbuf_1 _21219_ (.A(_05371_),
    .X(_01221_));
 sky130_fd_sc_hd__o211a_1 _21220_ (.A1(_05140_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05349_),
    .X(_05372_));
 sky130_fd_sc_hd__mux2_1 _21221_ (.A0(_05372_),
    .A1(net2464),
    .S(_05366_),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _21222_ (.A(_05373_),
    .X(_01222_));
 sky130_fd_sc_hd__o211a_1 _21223_ (.A1(_05143_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05352_),
    .X(_05374_));
 sky130_fd_sc_hd__mux2_1 _21224_ (.A0(_05374_),
    .A1(net3188),
    .S(_05366_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _21225_ (.A(_05375_),
    .X(_01223_));
 sky130_fd_sc_hd__o211a_1 _21226_ (.A1(_05146_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05355_),
    .X(_05376_));
 sky130_fd_sc_hd__mux2_1 _21227_ (.A0(_05376_),
    .A1(net3438),
    .S(_05366_),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _21228_ (.A(_05377_),
    .X(_01224_));
 sky130_fd_sc_hd__o211a_1 _21229_ (.A1(_05149_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05358_),
    .X(_05378_));
 sky130_fd_sc_hd__mux2_1 _21230_ (.A0(_05378_),
    .A1(net2990),
    .S(_05366_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _21231_ (.A(_05379_),
    .X(_01225_));
 sky130_fd_sc_hd__o211a_1 _21232_ (.A1(_05152_),
    .A2(_05338_),
    .B1(_05364_),
    .C1(_05361_),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _21233_ (.A0(_05380_),
    .A1(net3309),
    .S(_05366_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _21234_ (.A(_05381_),
    .X(_01226_));
 sky130_fd_sc_hd__o211a_1 _21235_ (.A1(_05059_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05340_),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_1 _21236_ (.A0(_05382_),
    .A1(net3289),
    .S(_05366_),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _21237_ (.A(_05383_),
    .X(_01227_));
 sky130_fd_sc_hd__o211a_1 _21238_ (.A1(_05063_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05343_),
    .X(_05384_));
 sky130_fd_sc_hd__mux2_1 _21239_ (.A0(_05384_),
    .A1(net3578),
    .S(_05366_),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _21240_ (.A(_05385_),
    .X(_01228_));
 sky130_fd_sc_hd__o211a_1 _21241_ (.A1(_05066_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05346_),
    .X(_05386_));
 sky130_fd_sc_hd__mux2_1 _21242_ (.A0(_05386_),
    .A1(net2661),
    .S(_05366_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _21243_ (.A(_05387_),
    .X(_01229_));
 sky130_fd_sc_hd__o211a_1 _21244_ (.A1(_05069_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05349_),
    .X(_05388_));
 sky130_fd_sc_hd__mux2_1 _21245_ (.A0(_05388_),
    .A1(net3388),
    .S(_05366_),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _21246_ (.A(_05389_),
    .X(_01230_));
 sky130_fd_sc_hd__o211a_1 _21247_ (.A1(_05072_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05352_),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _21248_ (.A0(_05390_),
    .A1(net2595),
    .S(_05366_),
    .X(_05391_));
 sky130_fd_sc_hd__clkbuf_1 _21249_ (.A(_05391_),
    .X(_01231_));
 sky130_fd_sc_hd__o211a_1 _21250_ (.A1(_05075_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05355_),
    .X(_05392_));
 sky130_fd_sc_hd__mux2_1 _21251_ (.A0(_05392_),
    .A1(net2688),
    .S(_05366_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _21252_ (.A(_05393_),
    .X(_01232_));
 sky130_fd_sc_hd__o211a_1 _21253_ (.A1(_05078_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05358_),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _21254_ (.A0(_05394_),
    .A1(net2306),
    .S(_05366_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _21255_ (.A(_05395_),
    .X(_01233_));
 sky130_fd_sc_hd__o211a_1 _21256_ (.A1(_05081_),
    .A2(_05339_),
    .B1(_05364_),
    .C1(_05361_),
    .X(_05396_));
 sky130_fd_sc_hd__mux2_1 _21257_ (.A0(_05396_),
    .A1(net2868),
    .S(_05366_),
    .X(_05397_));
 sky130_fd_sc_hd__clkbuf_1 _21258_ (.A(_05397_),
    .X(_01234_));
 sky130_fd_sc_hd__nand2_1 _21259_ (.A(_05319_),
    .B(_04183_),
    .Y(_05398_));
 sky130_fd_sc_hd__inv_2 _21260_ (.A(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__o21ai_4 _21261_ (.A1(_04332_),
    .A2(_05399_),
    .B1(_04776_),
    .Y(_05400_));
 sky130_fd_sc_hd__mux2_1 _21262_ (.A0(_05318_),
    .A1(net3270),
    .S(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _21263_ (.A(_05401_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _21264_ (.A0(_05324_),
    .A1(net3069),
    .S(_05400_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _21265_ (.A(_05402_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _21266_ (.A0(_05326_),
    .A1(net3649),
    .S(_05400_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _21267_ (.A(_05403_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _21268_ (.A0(_05328_),
    .A1(net2547),
    .S(_05400_),
    .X(_05404_));
 sky130_fd_sc_hd__clkbuf_1 _21269_ (.A(_05404_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _21270_ (.A0(_05330_),
    .A1(net3242),
    .S(_05400_),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_1 _21271_ (.A(_05405_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _21272_ (.A0(_05332_),
    .A1(net2566),
    .S(_05400_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _21273_ (.A(_05406_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _21274_ (.A0(_05334_),
    .A1(net3645),
    .S(_05400_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _21275_ (.A(_05407_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _21276_ (.A0(_05336_),
    .A1(net3320),
    .S(_05400_),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _21277_ (.A(_05408_),
    .X(_01242_));
 sky130_fd_sc_hd__buf_4 _21278_ (.A(_05400_),
    .X(_05409_));
 sky130_fd_sc_hd__buf_4 _21279_ (.A(_05399_),
    .X(_05410_));
 sky130_fd_sc_hd__buf_4 _21280_ (.A(_05399_),
    .X(_05411_));
 sky130_fd_sc_hd__nor2_1 _21281_ (.A(_02854_),
    .B(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__a211o_1 _21282_ (.A1(_02852_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_4 _21283_ (.A(_05400_),
    .X(_05414_));
 sky130_fd_sc_hd__nand2_1 _21284_ (.A(_05414_),
    .B(net552),
    .Y(_05415_));
 sky130_fd_sc_hd__o21ai_1 _21285_ (.A1(_05409_),
    .A2(_05413_),
    .B1(net553),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _21286_ (.A(_02863_),
    .B(_05411_),
    .Y(_05416_));
 sky130_fd_sc_hd__a211o_1 _21287_ (.A1(_02862_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__nand2_1 _21288_ (.A(_05414_),
    .B(net1987),
    .Y(_05418_));
 sky130_fd_sc_hd__o21ai_1 _21289_ (.A1(_05409_),
    .A2(_05417_),
    .B1(_05418_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _21290_ (.A(_02870_),
    .B(_05411_),
    .Y(_05419_));
 sky130_fd_sc_hd__a211o_1 _21291_ (.A1(_02869_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__nand2_1 _21292_ (.A(_05414_),
    .B(net512),
    .Y(_05421_));
 sky130_fd_sc_hd__o21ai_1 _21293_ (.A1(_05409_),
    .A2(_05420_),
    .B1(net513),
    .Y(_01245_));
 sky130_fd_sc_hd__nor2_1 _21294_ (.A(_02877_),
    .B(_05411_),
    .Y(_05422_));
 sky130_fd_sc_hd__a211o_1 _21295_ (.A1(_02876_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__nand2_1 _21296_ (.A(_05414_),
    .B(net536),
    .Y(_05424_));
 sky130_fd_sc_hd__o21ai_1 _21297_ (.A1(_05409_),
    .A2(_05423_),
    .B1(net537),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _21298_ (.A(_02884_),
    .B(_05411_),
    .Y(_05425_));
 sky130_fd_sc_hd__a211o_1 _21299_ (.A1(_02883_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__nand2_1 _21300_ (.A(_05414_),
    .B(net572),
    .Y(_05427_));
 sky130_fd_sc_hd__o21ai_1 _21301_ (.A1(_05409_),
    .A2(_05426_),
    .B1(net573),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _21302_ (.A(_02891_),
    .B(_05411_),
    .Y(_05428_));
 sky130_fd_sc_hd__a211o_1 _21303_ (.A1(_02890_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__nand2_1 _21304_ (.A(_05414_),
    .B(net1979),
    .Y(_05430_));
 sky130_fd_sc_hd__o21ai_1 _21305_ (.A1(_05409_),
    .A2(_05429_),
    .B1(_05430_),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _21306_ (.A(_02898_),
    .B(_05411_),
    .Y(_05431_));
 sky130_fd_sc_hd__a211o_1 _21307_ (.A1(_02897_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__nand2_1 _21308_ (.A(_05414_),
    .B(net1808),
    .Y(_05433_));
 sky130_fd_sc_hd__o21ai_1 _21309_ (.A1(_05409_),
    .A2(_05432_),
    .B1(net1809),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_1 _21310_ (.A(_02905_),
    .B(_05411_),
    .Y(_05434_));
 sky130_fd_sc_hd__a211o_1 _21311_ (.A1(_02904_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__nand2_1 _21312_ (.A(_05414_),
    .B(net472),
    .Y(_05436_));
 sky130_fd_sc_hd__o21ai_1 _21313_ (.A1(_05409_),
    .A2(_05435_),
    .B1(net473),
    .Y(_01250_));
 sky130_fd_sc_hd__buf_4 _21314_ (.A(_05400_),
    .X(_05437_));
 sky130_fd_sc_hd__a211o_1 _21315_ (.A1(_02912_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05412_),
    .X(_05438_));
 sky130_fd_sc_hd__nand2_1 _21316_ (.A(_05414_),
    .B(net1488),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_1 _21317_ (.A1(_05437_),
    .A2(_05438_),
    .B1(net1489),
    .Y(_01251_));
 sky130_fd_sc_hd__a211o_1 _21318_ (.A1(_02917_),
    .A2(_05410_),
    .B1(_05305_),
    .C1(_05416_),
    .X(_05440_));
 sky130_fd_sc_hd__nand2_1 _21319_ (.A(_05414_),
    .B(net1494),
    .Y(_05441_));
 sky130_fd_sc_hd__o21ai_1 _21320_ (.A1(_05437_),
    .A2(_05440_),
    .B1(net1495),
    .Y(_01252_));
 sky130_fd_sc_hd__buf_4 _21321_ (.A(_04598_),
    .X(_05442_));
 sky130_fd_sc_hd__a211o_1 _21322_ (.A1(_02922_),
    .A2(_05410_),
    .B1(_05442_),
    .C1(_05419_),
    .X(_05443_));
 sky130_fd_sc_hd__nand2_1 _21323_ (.A(_05414_),
    .B(net1114),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_1 _21324_ (.A1(_05437_),
    .A2(_05443_),
    .B1(net1115),
    .Y(_01253_));
 sky130_fd_sc_hd__a211o_1 _21325_ (.A1(_02928_),
    .A2(_05410_),
    .B1(_05442_),
    .C1(_05422_),
    .X(_05445_));
 sky130_fd_sc_hd__nand2_1 _21326_ (.A(_05414_),
    .B(net1290),
    .Y(_05446_));
 sky130_fd_sc_hd__o21ai_1 _21327_ (.A1(_05437_),
    .A2(_05445_),
    .B1(net1291),
    .Y(_01254_));
 sky130_fd_sc_hd__a211o_1 _21328_ (.A1(_02933_),
    .A2(_05410_),
    .B1(_05442_),
    .C1(_05425_),
    .X(_05447_));
 sky130_fd_sc_hd__nand2_1 _21329_ (.A(_05414_),
    .B(net856),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_1 _21330_ (.A1(_05437_),
    .A2(_05447_),
    .B1(net857),
    .Y(_01255_));
 sky130_fd_sc_hd__a211o_1 _21331_ (.A1(_02938_),
    .A2(_05410_),
    .B1(_05442_),
    .C1(_05428_),
    .X(_05449_));
 sky130_fd_sc_hd__nand2_1 _21332_ (.A(_05414_),
    .B(net858),
    .Y(_05450_));
 sky130_fd_sc_hd__o21ai_1 _21333_ (.A1(_05437_),
    .A2(_05449_),
    .B1(net859),
    .Y(_01256_));
 sky130_fd_sc_hd__a211o_1 _21334_ (.A1(_02943_),
    .A2(_05410_),
    .B1(_05442_),
    .C1(_05431_),
    .X(_05451_));
 sky130_fd_sc_hd__nand2_1 _21335_ (.A(_05414_),
    .B(net1670),
    .Y(_05452_));
 sky130_fd_sc_hd__o21ai_1 _21336_ (.A1(_05437_),
    .A2(_05451_),
    .B1(net1671),
    .Y(_01257_));
 sky130_fd_sc_hd__a211o_1 _21337_ (.A1(_02948_),
    .A2(_05410_),
    .B1(_05442_),
    .C1(_05434_),
    .X(_05453_));
 sky130_fd_sc_hd__nand2_1 _21338_ (.A(_05414_),
    .B(net1450),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ai_1 _21339_ (.A1(_05437_),
    .A2(_05453_),
    .B1(net1451),
    .Y(_01258_));
 sky130_fd_sc_hd__a211o_1 _21340_ (.A1(_02952_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05412_),
    .X(_05455_));
 sky130_fd_sc_hd__nand2_1 _21341_ (.A(_05409_),
    .B(net1402),
    .Y(_05456_));
 sky130_fd_sc_hd__o21ai_1 _21342_ (.A1(_05437_),
    .A2(_05455_),
    .B1(net1403),
    .Y(_01259_));
 sky130_fd_sc_hd__a211o_1 _21343_ (.A1(_02956_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05416_),
    .X(_05457_));
 sky130_fd_sc_hd__nand2_1 _21344_ (.A(_05409_),
    .B(net1326),
    .Y(_05458_));
 sky130_fd_sc_hd__o21ai_1 _21345_ (.A1(_05437_),
    .A2(_05457_),
    .B1(net1327),
    .Y(_01260_));
 sky130_fd_sc_hd__a211o_1 _21346_ (.A1(_02960_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05419_),
    .X(_05459_));
 sky130_fd_sc_hd__nand2_1 _21347_ (.A(_05409_),
    .B(net1830),
    .Y(_05460_));
 sky130_fd_sc_hd__o21ai_1 _21348_ (.A1(_05437_),
    .A2(_05459_),
    .B1(net1831),
    .Y(_01261_));
 sky130_fd_sc_hd__a211o_1 _21349_ (.A1(_02964_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05422_),
    .X(_05461_));
 sky130_fd_sc_hd__nand2_1 _21350_ (.A(_05409_),
    .B(net1280),
    .Y(_05462_));
 sky130_fd_sc_hd__o21ai_1 _21351_ (.A1(_05437_),
    .A2(_05461_),
    .B1(net1281),
    .Y(_01262_));
 sky130_fd_sc_hd__a211o_1 _21352_ (.A1(_02968_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05425_),
    .X(_05463_));
 sky130_fd_sc_hd__nand2_1 _21353_ (.A(_05409_),
    .B(net1250),
    .Y(_05464_));
 sky130_fd_sc_hd__o21ai_1 _21354_ (.A1(_05437_),
    .A2(_05463_),
    .B1(net1251),
    .Y(_01263_));
 sky130_fd_sc_hd__a211o_1 _21355_ (.A1(_02972_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05428_),
    .X(_05465_));
 sky130_fd_sc_hd__nand2_1 _21356_ (.A(_05409_),
    .B(net1756),
    .Y(_05466_));
 sky130_fd_sc_hd__o21ai_1 _21357_ (.A1(_05437_),
    .A2(_05465_),
    .B1(net1757),
    .Y(_01264_));
 sky130_fd_sc_hd__a211o_1 _21358_ (.A1(_02976_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05431_),
    .X(_05467_));
 sky130_fd_sc_hd__nand2_1 _21359_ (.A(_05409_),
    .B(net1268),
    .Y(_05468_));
 sky130_fd_sc_hd__o21ai_1 _21360_ (.A1(_05437_),
    .A2(_05467_),
    .B1(net1269),
    .Y(_01265_));
 sky130_fd_sc_hd__a211o_1 _21361_ (.A1(_02980_),
    .A2(_05411_),
    .B1(_05442_),
    .C1(_05434_),
    .X(_05469_));
 sky130_fd_sc_hd__nand2_1 _21362_ (.A(_05409_),
    .B(net1082),
    .Y(_05470_));
 sky130_fd_sc_hd__o21ai_1 _21363_ (.A1(_05437_),
    .A2(_05469_),
    .B1(net1083),
    .Y(_01266_));
 sky130_fd_sc_hd__buf_12 _21364_ (.A(_12289_),
    .X(_05471_));
 sky130_fd_sc_hd__nand2_1 _21365_ (.A(_05319_),
    .B(_04257_),
    .Y(_05472_));
 sky130_fd_sc_hd__inv_2 _21366_ (.A(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21ai_4 _21367_ (.A1(_05471_),
    .A2(_05473_),
    .B1(_04776_),
    .Y(_05474_));
 sky130_fd_sc_hd__mux2_1 _21368_ (.A0(_05318_),
    .A1(net3293),
    .S(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__clkbuf_1 _21369_ (.A(_05475_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _21370_ (.A0(_05324_),
    .A1(net3545),
    .S(_05474_),
    .X(_05476_));
 sky130_fd_sc_hd__clkbuf_1 _21371_ (.A(_05476_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _21372_ (.A0(_05326_),
    .A1(net2903),
    .S(_05474_),
    .X(_05477_));
 sky130_fd_sc_hd__clkbuf_1 _21373_ (.A(_05477_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _21374_ (.A0(_05328_),
    .A1(net3034),
    .S(_05474_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_1 _21375_ (.A(_05478_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _21376_ (.A0(_05330_),
    .A1(net3489),
    .S(_05474_),
    .X(_05479_));
 sky130_fd_sc_hd__clkbuf_1 _21377_ (.A(_05479_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _21378_ (.A0(_05332_),
    .A1(net3424),
    .S(_05474_),
    .X(_05480_));
 sky130_fd_sc_hd__clkbuf_1 _21379_ (.A(_05480_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _21380_ (.A0(_05334_),
    .A1(net3060),
    .S(_05474_),
    .X(_05481_));
 sky130_fd_sc_hd__clkbuf_1 _21381_ (.A(_05481_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _21382_ (.A0(_05336_),
    .A1(net2980),
    .S(_05474_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _21383_ (.A(_05482_),
    .X(_01274_));
 sky130_fd_sc_hd__buf_4 _21384_ (.A(_05474_),
    .X(_05483_));
 sky130_fd_sc_hd__clkbuf_16 _21385_ (.A(_02851_),
    .X(_05484_));
 sky130_fd_sc_hd__buf_4 _21386_ (.A(_05473_),
    .X(_05485_));
 sky130_fd_sc_hd__buf_4 _21387_ (.A(_05473_),
    .X(_05486_));
 sky130_fd_sc_hd__nor2_1 _21388_ (.A(_02854_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__a211o_1 _21389_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05442_),
    .C1(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__buf_4 _21390_ (.A(_05474_),
    .X(_05489_));
 sky130_fd_sc_hd__nand2_1 _21391_ (.A(_05489_),
    .B(net726),
    .Y(_05490_));
 sky130_fd_sc_hd__o21ai_1 _21392_ (.A1(_05483_),
    .A2(_05488_),
    .B1(net727),
    .Y(_01275_));
 sky130_fd_sc_hd__clkbuf_16 _21393_ (.A(_02861_),
    .X(_05491_));
 sky130_fd_sc_hd__nor2_1 _21394_ (.A(_02863_),
    .B(_05486_),
    .Y(_05492_));
 sky130_fd_sc_hd__a211o_1 _21395_ (.A1(_05491_),
    .A2(_05485_),
    .B1(_05442_),
    .C1(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__nand2_1 _21396_ (.A(_05489_),
    .B(net922),
    .Y(_05494_));
 sky130_fd_sc_hd__o21ai_1 _21397_ (.A1(_05483_),
    .A2(_05493_),
    .B1(net923),
    .Y(_01276_));
 sky130_fd_sc_hd__clkbuf_16 _21398_ (.A(_02868_),
    .X(_05495_));
 sky130_fd_sc_hd__buf_4 _21399_ (.A(_04598_),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_1 _21400_ (.A(_02870_),
    .B(_05486_),
    .Y(_05497_));
 sky130_fd_sc_hd__a211o_1 _21401_ (.A1(_05495_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__nand2_1 _21402_ (.A(_05489_),
    .B(net764),
    .Y(_05499_));
 sky130_fd_sc_hd__o21ai_1 _21403_ (.A1(_05483_),
    .A2(_05498_),
    .B1(net765),
    .Y(_01277_));
 sky130_fd_sc_hd__clkbuf_16 _21404_ (.A(_02875_),
    .X(_05500_));
 sky130_fd_sc_hd__nor2_1 _21405_ (.A(_02877_),
    .B(_05486_),
    .Y(_05501_));
 sky130_fd_sc_hd__a211o_1 _21406_ (.A1(_05500_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__nand2_1 _21407_ (.A(_05489_),
    .B(net712),
    .Y(_05503_));
 sky130_fd_sc_hd__o21ai_1 _21408_ (.A1(_05483_),
    .A2(_05502_),
    .B1(net713),
    .Y(_01278_));
 sky130_fd_sc_hd__clkbuf_16 _21409_ (.A(_02882_),
    .X(_05504_));
 sky130_fd_sc_hd__nor2_1 _21410_ (.A(_02884_),
    .B(_05486_),
    .Y(_05505_));
 sky130_fd_sc_hd__a211o_1 _21411_ (.A1(_05504_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__nand2_1 _21412_ (.A(_05489_),
    .B(net1190),
    .Y(_05507_));
 sky130_fd_sc_hd__o21ai_1 _21413_ (.A1(_05483_),
    .A2(_05506_),
    .B1(net1191),
    .Y(_01279_));
 sky130_fd_sc_hd__clkbuf_16 _21414_ (.A(_02889_),
    .X(_05508_));
 sky130_fd_sc_hd__nor2_1 _21415_ (.A(_02891_),
    .B(_05486_),
    .Y(_05509_));
 sky130_fd_sc_hd__a211o_1 _21416_ (.A1(_05508_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__nand2_1 _21417_ (.A(_05489_),
    .B(net988),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_1 _21418_ (.A1(_05483_),
    .A2(_05510_),
    .B1(net989),
    .Y(_01280_));
 sky130_fd_sc_hd__clkbuf_16 _21419_ (.A(_02896_),
    .X(_05512_));
 sky130_fd_sc_hd__nor2_1 _21420_ (.A(_02898_),
    .B(_05486_),
    .Y(_05513_));
 sky130_fd_sc_hd__a211o_1 _21421_ (.A1(_05512_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__nand2_1 _21422_ (.A(_05489_),
    .B(net876),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_1 _21423_ (.A1(_05483_),
    .A2(_05514_),
    .B1(net877),
    .Y(_01281_));
 sky130_fd_sc_hd__clkbuf_16 _21424_ (.A(_02903_),
    .X(_05516_));
 sky130_fd_sc_hd__nor2_1 _21425_ (.A(_02905_),
    .B(_05486_),
    .Y(_05517_));
 sky130_fd_sc_hd__a211o_1 _21426_ (.A1(_05516_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__nand2_1 _21427_ (.A(_05489_),
    .B(net668),
    .Y(_05519_));
 sky130_fd_sc_hd__o21ai_1 _21428_ (.A1(_05483_),
    .A2(_05518_),
    .B1(net669),
    .Y(_01282_));
 sky130_fd_sc_hd__buf_4 _21429_ (.A(_05474_),
    .X(_05520_));
 sky130_fd_sc_hd__buf_12 _21430_ (.A(_02911_),
    .X(_05521_));
 sky130_fd_sc_hd__a211o_1 _21431_ (.A1(_05521_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05487_),
    .X(_05522_));
 sky130_fd_sc_hd__nand2_1 _21432_ (.A(_05489_),
    .B(net1012),
    .Y(_05523_));
 sky130_fd_sc_hd__o21ai_1 _21433_ (.A1(_05520_),
    .A2(_05522_),
    .B1(net1013),
    .Y(_01283_));
 sky130_fd_sc_hd__clkbuf_16 _21434_ (.A(_02916_),
    .X(_05524_));
 sky130_fd_sc_hd__a211o_1 _21435_ (.A1(_05524_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05492_),
    .X(_05525_));
 sky130_fd_sc_hd__nand2_1 _21436_ (.A(_05489_),
    .B(net1528),
    .Y(_05526_));
 sky130_fd_sc_hd__o21ai_1 _21437_ (.A1(_05520_),
    .A2(_05525_),
    .B1(net1529),
    .Y(_01284_));
 sky130_fd_sc_hd__clkbuf_16 _21438_ (.A(_02921_),
    .X(_05527_));
 sky130_fd_sc_hd__a211o_1 _21439_ (.A1(_05527_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05497_),
    .X(_05528_));
 sky130_fd_sc_hd__nand2_1 _21440_ (.A(_05489_),
    .B(net1873),
    .Y(_05529_));
 sky130_fd_sc_hd__o21ai_1 _21441_ (.A1(_05520_),
    .A2(_05528_),
    .B1(net1874),
    .Y(_01285_));
 sky130_fd_sc_hd__buf_12 _21442_ (.A(_02927_),
    .X(_05530_));
 sky130_fd_sc_hd__a211o_1 _21443_ (.A1(_05530_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05501_),
    .X(_05531_));
 sky130_fd_sc_hd__nand2_1 _21444_ (.A(_05489_),
    .B(net710),
    .Y(_05532_));
 sky130_fd_sc_hd__o21ai_1 _21445_ (.A1(_05520_),
    .A2(_05531_),
    .B1(net711),
    .Y(_01286_));
 sky130_fd_sc_hd__clkbuf_16 _21446_ (.A(_02932_),
    .X(_05533_));
 sky130_fd_sc_hd__a211o_1 _21447_ (.A1(_05533_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05505_),
    .X(_05534_));
 sky130_fd_sc_hd__nand2_1 _21448_ (.A(_05489_),
    .B(net1024),
    .Y(_05535_));
 sky130_fd_sc_hd__o21ai_1 _21449_ (.A1(_05520_),
    .A2(_05534_),
    .B1(net1025),
    .Y(_01287_));
 sky130_fd_sc_hd__clkbuf_16 _21450_ (.A(_02937_),
    .X(_05536_));
 sky130_fd_sc_hd__a211o_1 _21451_ (.A1(_05536_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05509_),
    .X(_05537_));
 sky130_fd_sc_hd__nand2_1 _21452_ (.A(_05489_),
    .B(net932),
    .Y(_05538_));
 sky130_fd_sc_hd__o21ai_1 _21453_ (.A1(_05520_),
    .A2(_05537_),
    .B1(net933),
    .Y(_01288_));
 sky130_fd_sc_hd__clkbuf_16 _21454_ (.A(_02942_),
    .X(_05539_));
 sky130_fd_sc_hd__a211o_1 _21455_ (.A1(_05539_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05513_),
    .X(_05540_));
 sky130_fd_sc_hd__nand2_1 _21456_ (.A(_05489_),
    .B(net1624),
    .Y(_05541_));
 sky130_fd_sc_hd__o21ai_1 _21457_ (.A1(_05520_),
    .A2(_05540_),
    .B1(net1625),
    .Y(_01289_));
 sky130_fd_sc_hd__clkbuf_16 _21458_ (.A(_02947_),
    .X(_05542_));
 sky130_fd_sc_hd__a211o_1 _21459_ (.A1(_05542_),
    .A2(_05485_),
    .B1(_05496_),
    .C1(_05517_),
    .X(_05543_));
 sky130_fd_sc_hd__nand2_1 _21460_ (.A(_05489_),
    .B(net1762),
    .Y(_05544_));
 sky130_fd_sc_hd__o21ai_1 _21461_ (.A1(_05520_),
    .A2(_05543_),
    .B1(net1763),
    .Y(_01290_));
 sky130_fd_sc_hd__clkbuf_16 _21462_ (.A(_02951_),
    .X(_05545_));
 sky130_fd_sc_hd__a211o_1 _21463_ (.A1(_05545_),
    .A2(_05486_),
    .B1(_05496_),
    .C1(_05487_),
    .X(_05546_));
 sky130_fd_sc_hd__nand2_1 _21464_ (.A(_05483_),
    .B(net692),
    .Y(_05547_));
 sky130_fd_sc_hd__o21ai_1 _21465_ (.A1(_05520_),
    .A2(_05546_),
    .B1(net693),
    .Y(_01291_));
 sky130_fd_sc_hd__buf_12 _21466_ (.A(_02955_),
    .X(_05548_));
 sky130_fd_sc_hd__a211o_1 _21467_ (.A1(_05548_),
    .A2(_05486_),
    .B1(_05496_),
    .C1(_05492_),
    .X(_05549_));
 sky130_fd_sc_hd__nand2_1 _21468_ (.A(_05483_),
    .B(net782),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_1 _21469_ (.A1(_05520_),
    .A2(_05549_),
    .B1(net783),
    .Y(_01292_));
 sky130_fd_sc_hd__clkbuf_16 _21470_ (.A(_02959_),
    .X(_05551_));
 sky130_fd_sc_hd__buf_4 _21471_ (.A(_04598_),
    .X(_05552_));
 sky130_fd_sc_hd__a211o_1 _21472_ (.A1(_05551_),
    .A2(_05486_),
    .B1(_05552_),
    .C1(_05497_),
    .X(_05553_));
 sky130_fd_sc_hd__nand2_1 _21473_ (.A(_05483_),
    .B(net1824),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_1 _21474_ (.A1(_05520_),
    .A2(_05553_),
    .B1(net1825),
    .Y(_01293_));
 sky130_fd_sc_hd__buf_12 _21475_ (.A(_02963_),
    .X(_05555_));
 sky130_fd_sc_hd__a211o_1 _21476_ (.A1(_05555_),
    .A2(_05486_),
    .B1(_05552_),
    .C1(_05501_),
    .X(_05556_));
 sky130_fd_sc_hd__nand2_1 _21477_ (.A(_05483_),
    .B(net1084),
    .Y(_05557_));
 sky130_fd_sc_hd__o21ai_1 _21478_ (.A1(_05520_),
    .A2(_05556_),
    .B1(net1085),
    .Y(_01294_));
 sky130_fd_sc_hd__clkbuf_16 _21479_ (.A(_02967_),
    .X(_05558_));
 sky130_fd_sc_hd__a211o_1 _21480_ (.A1(_05558_),
    .A2(_05486_),
    .B1(_05552_),
    .C1(_05505_),
    .X(_05559_));
 sky130_fd_sc_hd__nand2_1 _21481_ (.A(_05483_),
    .B(net1786),
    .Y(_05560_));
 sky130_fd_sc_hd__o21ai_1 _21482_ (.A1(_05520_),
    .A2(_05559_),
    .B1(net1787),
    .Y(_01295_));
 sky130_fd_sc_hd__clkbuf_16 _21483_ (.A(_02971_),
    .X(_05561_));
 sky130_fd_sc_hd__a211o_1 _21484_ (.A1(_05561_),
    .A2(_05486_),
    .B1(_05552_),
    .C1(_05509_),
    .X(_05562_));
 sky130_fd_sc_hd__nand2_1 _21485_ (.A(_05483_),
    .B(net1752),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ai_1 _21486_ (.A1(_05520_),
    .A2(_05562_),
    .B1(net1753),
    .Y(_01296_));
 sky130_fd_sc_hd__clkbuf_16 _21487_ (.A(_02975_),
    .X(_05564_));
 sky130_fd_sc_hd__a211o_1 _21488_ (.A1(_05564_),
    .A2(_05486_),
    .B1(_05552_),
    .C1(_05513_),
    .X(_05565_));
 sky130_fd_sc_hd__nand2_1 _21489_ (.A(_05483_),
    .B(net1380),
    .Y(_05566_));
 sky130_fd_sc_hd__o21ai_1 _21490_ (.A1(_05520_),
    .A2(_05565_),
    .B1(net1381),
    .Y(_01297_));
 sky130_fd_sc_hd__buf_12 _21491_ (.A(_02979_),
    .X(_05567_));
 sky130_fd_sc_hd__a211o_1 _21492_ (.A1(_05567_),
    .A2(_05486_),
    .B1(_05552_),
    .C1(_05517_),
    .X(_05568_));
 sky130_fd_sc_hd__nand2_1 _21493_ (.A(_05483_),
    .B(net1136),
    .Y(_05569_));
 sky130_fd_sc_hd__o21ai_1 _21494_ (.A1(_05520_),
    .A2(_05568_),
    .B1(net1137),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _21495_ (.A(_05319_),
    .B(_04333_),
    .Y(_05570_));
 sky130_fd_sc_hd__inv_2 _21496_ (.A(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21ai_4 _21497_ (.A1(_05471_),
    .A2(_05571_),
    .B1(_04776_),
    .Y(_05572_));
 sky130_fd_sc_hd__mux2_1 _21498_ (.A0(_05318_),
    .A1(net2789),
    .S(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _21499_ (.A(_05573_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _21500_ (.A0(_05324_),
    .A1(net2521),
    .S(_05572_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _21501_ (.A(_05574_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _21502_ (.A0(_05326_),
    .A1(net3297),
    .S(_05572_),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_1 _21503_ (.A(_05575_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _21504_ (.A0(_05328_),
    .A1(net2289),
    .S(_05572_),
    .X(_05576_));
 sky130_fd_sc_hd__clkbuf_1 _21505_ (.A(_05576_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _21506_ (.A0(_05330_),
    .A1(net2803),
    .S(_05572_),
    .X(_05577_));
 sky130_fd_sc_hd__clkbuf_1 _21507_ (.A(_05577_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _21508_ (.A0(_05332_),
    .A1(net3433),
    .S(_05572_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_1 _21509_ (.A(_05578_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _21510_ (.A0(_05334_),
    .A1(net2981),
    .S(_05572_),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_1 _21511_ (.A(_05579_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _21512_ (.A0(_05336_),
    .A1(net3166),
    .S(_05572_),
    .X(_05580_));
 sky130_fd_sc_hd__clkbuf_1 _21513_ (.A(_05580_),
    .X(_01306_));
 sky130_fd_sc_hd__buf_4 _21514_ (.A(_05572_),
    .X(_05581_));
 sky130_fd_sc_hd__buf_4 _21515_ (.A(_05571_),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_16 _21516_ (.A(_12183_),
    .X(_05583_));
 sky130_fd_sc_hd__buf_4 _21517_ (.A(_05571_),
    .X(_05584_));
 sky130_fd_sc_hd__nor2_1 _21518_ (.A(_05583_),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a211o_1 _21519_ (.A1(_05484_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_4 _21520_ (.A(_05572_),
    .X(_05587_));
 sky130_fd_sc_hd__nand2_1 _21521_ (.A(_05587_),
    .B(net1260),
    .Y(_05588_));
 sky130_fd_sc_hd__o21ai_1 _21522_ (.A1(_05581_),
    .A2(_05586_),
    .B1(net1261),
    .Y(_01307_));
 sky130_fd_sc_hd__clkbuf_16 _21523_ (.A(_12196_),
    .X(_05589_));
 sky130_fd_sc_hd__nor2_1 _21524_ (.A(_05589_),
    .B(_05584_),
    .Y(_05590_));
 sky130_fd_sc_hd__a211o_1 _21525_ (.A1(_05491_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__nand2_1 _21526_ (.A(_05587_),
    .B(net1408),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ai_1 _21527_ (.A1(_05581_),
    .A2(_05591_),
    .B1(net1409),
    .Y(_01308_));
 sky130_fd_sc_hd__buf_12 _21528_ (.A(_12204_),
    .X(_05593_));
 sky130_fd_sc_hd__nor2_1 _21529_ (.A(_05593_),
    .B(_05584_),
    .Y(_05594_));
 sky130_fd_sc_hd__a211o_1 _21530_ (.A1(_05495_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__nand2_1 _21531_ (.A(_05587_),
    .B(net1428),
    .Y(_05596_));
 sky130_fd_sc_hd__o21ai_1 _21532_ (.A1(_05581_),
    .A2(_05595_),
    .B1(net1429),
    .Y(_01309_));
 sky130_fd_sc_hd__clkbuf_16 _21533_ (.A(_12212_),
    .X(_05597_));
 sky130_fd_sc_hd__nor2_1 _21534_ (.A(_05597_),
    .B(_05584_),
    .Y(_05598_));
 sky130_fd_sc_hd__a211o_1 _21535_ (.A1(_05500_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__nand2_1 _21536_ (.A(_05587_),
    .B(net680),
    .Y(_05600_));
 sky130_fd_sc_hd__o21ai_1 _21537_ (.A1(_05581_),
    .A2(_05599_),
    .B1(net681),
    .Y(_01310_));
 sky130_fd_sc_hd__clkbuf_16 _21538_ (.A(_12220_),
    .X(_05601_));
 sky130_fd_sc_hd__nor2_1 _21539_ (.A(_05601_),
    .B(_05584_),
    .Y(_05602_));
 sky130_fd_sc_hd__a211o_1 _21540_ (.A1(_05504_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__nand2_1 _21541_ (.A(_05587_),
    .B(net1066),
    .Y(_05604_));
 sky130_fd_sc_hd__o21ai_1 _21542_ (.A1(_05581_),
    .A2(_05603_),
    .B1(net1067),
    .Y(_01311_));
 sky130_fd_sc_hd__clkbuf_16 _21543_ (.A(_12228_),
    .X(_05605_));
 sky130_fd_sc_hd__nor2_1 _21544_ (.A(_05605_),
    .B(_05584_),
    .Y(_05606_));
 sky130_fd_sc_hd__a211o_1 _21545_ (.A1(_05508_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__nand2_1 _21546_ (.A(_05587_),
    .B(net1342),
    .Y(_05608_));
 sky130_fd_sc_hd__o21ai_1 _21547_ (.A1(_05581_),
    .A2(_05607_),
    .B1(net1343),
    .Y(_01312_));
 sky130_fd_sc_hd__buf_12 _21548_ (.A(_12236_),
    .X(_05609_));
 sky130_fd_sc_hd__nor2_1 _21549_ (.A(_05609_),
    .B(_05584_),
    .Y(_05610_));
 sky130_fd_sc_hd__a211o_1 _21550_ (.A1(_05512_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__nand2_1 _21551_ (.A(_05587_),
    .B(net522),
    .Y(_05612_));
 sky130_fd_sc_hd__o21ai_1 _21552_ (.A1(_05581_),
    .A2(_05611_),
    .B1(net523),
    .Y(_01313_));
 sky130_fd_sc_hd__clkbuf_16 _21553_ (.A(_12244_),
    .X(_05613_));
 sky130_fd_sc_hd__nor2_1 _21554_ (.A(_05613_),
    .B(_05584_),
    .Y(_05614_));
 sky130_fd_sc_hd__a211o_1 _21555_ (.A1(_05516_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__nand2_1 _21556_ (.A(_05587_),
    .B(net498),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_1 _21557_ (.A1(_05581_),
    .A2(_05615_),
    .B1(net499),
    .Y(_01314_));
 sky130_fd_sc_hd__buf_4 _21558_ (.A(_05572_),
    .X(_05617_));
 sky130_fd_sc_hd__a211o_1 _21559_ (.A1(_05521_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05585_),
    .X(_05618_));
 sky130_fd_sc_hd__nand2_1 _21560_ (.A(_05587_),
    .B(net1622),
    .Y(_05619_));
 sky130_fd_sc_hd__o21ai_1 _21561_ (.A1(_05617_),
    .A2(_05618_),
    .B1(net1623),
    .Y(_01315_));
 sky130_fd_sc_hd__a211o_1 _21562_ (.A1(_05524_),
    .A2(_05582_),
    .B1(_05552_),
    .C1(_05590_),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_1 _21563_ (.A(_05587_),
    .B(net966),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_1 _21564_ (.A1(_05617_),
    .A2(_05620_),
    .B1(net967),
    .Y(_01316_));
 sky130_fd_sc_hd__buf_4 _21565_ (.A(_04598_),
    .X(_05622_));
 sky130_fd_sc_hd__a211o_1 _21566_ (.A1(_05527_),
    .A2(_05582_),
    .B1(_05622_),
    .C1(_05594_),
    .X(_05623_));
 sky130_fd_sc_hd__nand2_1 _21567_ (.A(_05587_),
    .B(net924),
    .Y(_05624_));
 sky130_fd_sc_hd__o21ai_1 _21568_ (.A1(_05617_),
    .A2(_05623_),
    .B1(net925),
    .Y(_01317_));
 sky130_fd_sc_hd__a211o_1 _21569_ (.A1(_05530_),
    .A2(_05582_),
    .B1(_05622_),
    .C1(_05598_),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _21570_ (.A(_05587_),
    .B(net1098),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_1 _21571_ (.A1(_05617_),
    .A2(_05625_),
    .B1(net1099),
    .Y(_01318_));
 sky130_fd_sc_hd__a211o_1 _21572_ (.A1(_05533_),
    .A2(_05582_),
    .B1(_05622_),
    .C1(_05602_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _21573_ (.A(_05587_),
    .B(net1680),
    .Y(_05628_));
 sky130_fd_sc_hd__o21ai_1 _21574_ (.A1(_05617_),
    .A2(_05627_),
    .B1(net1681),
    .Y(_01319_));
 sky130_fd_sc_hd__a211o_1 _21575_ (.A1(_05536_),
    .A2(_05582_),
    .B1(_05622_),
    .C1(_05606_),
    .X(_05629_));
 sky130_fd_sc_hd__nand2_1 _21576_ (.A(_05587_),
    .B(net1346),
    .Y(_05630_));
 sky130_fd_sc_hd__o21ai_1 _21577_ (.A1(_05617_),
    .A2(_05629_),
    .B1(net1347),
    .Y(_01320_));
 sky130_fd_sc_hd__a211o_1 _21578_ (.A1(_05539_),
    .A2(_05582_),
    .B1(_05622_),
    .C1(_05610_),
    .X(_05631_));
 sky130_fd_sc_hd__nand2_1 _21579_ (.A(_05587_),
    .B(net1302),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_1 _21580_ (.A1(_05617_),
    .A2(_05631_),
    .B1(net1303),
    .Y(_01321_));
 sky130_fd_sc_hd__a211o_1 _21581_ (.A1(_05542_),
    .A2(_05582_),
    .B1(_05622_),
    .C1(_05614_),
    .X(_05633_));
 sky130_fd_sc_hd__nand2_1 _21582_ (.A(_05587_),
    .B(net866),
    .Y(_05634_));
 sky130_fd_sc_hd__o21ai_1 _21583_ (.A1(_05617_),
    .A2(_05633_),
    .B1(net867),
    .Y(_01322_));
 sky130_fd_sc_hd__a211o_1 _21584_ (.A1(_05545_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05585_),
    .X(_05635_));
 sky130_fd_sc_hd__nand2_1 _21585_ (.A(_05581_),
    .B(net1108),
    .Y(_05636_));
 sky130_fd_sc_hd__o21ai_1 _21586_ (.A1(_05617_),
    .A2(_05635_),
    .B1(net1109),
    .Y(_01323_));
 sky130_fd_sc_hd__a211o_1 _21587_ (.A1(_05548_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05590_),
    .X(_05637_));
 sky130_fd_sc_hd__nand2_1 _21588_ (.A(_05581_),
    .B(net1142),
    .Y(_05638_));
 sky130_fd_sc_hd__o21ai_1 _21589_ (.A1(_05617_),
    .A2(_05637_),
    .B1(net1143),
    .Y(_01324_));
 sky130_fd_sc_hd__a211o_1 _21590_ (.A1(_05551_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05594_),
    .X(_05639_));
 sky130_fd_sc_hd__nand2_1 _21591_ (.A(_05581_),
    .B(net918),
    .Y(_05640_));
 sky130_fd_sc_hd__o21ai_1 _21592_ (.A1(_05617_),
    .A2(_05639_),
    .B1(net919),
    .Y(_01325_));
 sky130_fd_sc_hd__a211o_1 _21593_ (.A1(_05555_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05598_),
    .X(_05641_));
 sky130_fd_sc_hd__nand2_1 _21594_ (.A(_05581_),
    .B(net1242),
    .Y(_05642_));
 sky130_fd_sc_hd__o21ai_1 _21595_ (.A1(_05617_),
    .A2(_05641_),
    .B1(net1243),
    .Y(_01326_));
 sky130_fd_sc_hd__a211o_1 _21596_ (.A1(_05558_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05602_),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_1 _21597_ (.A(_05581_),
    .B(net1730),
    .Y(_05644_));
 sky130_fd_sc_hd__o21ai_1 _21598_ (.A1(_05617_),
    .A2(_05643_),
    .B1(net1731),
    .Y(_01327_));
 sky130_fd_sc_hd__a211o_1 _21599_ (.A1(_05561_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05606_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _21600_ (.A(_05581_),
    .B(net826),
    .Y(_05646_));
 sky130_fd_sc_hd__o21ai_1 _21601_ (.A1(_05617_),
    .A2(_05645_),
    .B1(net827),
    .Y(_01328_));
 sky130_fd_sc_hd__a211o_1 _21602_ (.A1(_05564_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05610_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _21603_ (.A(_05581_),
    .B(net1230),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_1 _21604_ (.A1(_05617_),
    .A2(_05647_),
    .B1(net1231),
    .Y(_01329_));
 sky130_fd_sc_hd__a211o_1 _21605_ (.A1(_05567_),
    .A2(_05584_),
    .B1(_05622_),
    .C1(_05614_),
    .X(_05649_));
 sky130_fd_sc_hd__nand2_1 _21606_ (.A(_05581_),
    .B(net1480),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_1 _21607_ (.A1(_05617_),
    .A2(_05649_),
    .B1(net1481),
    .Y(_01330_));
 sky130_fd_sc_hd__and3_2 _21608_ (.A(_03207_),
    .B(\line_cache_idx[7] ),
    .C(_12303_),
    .X(_05651_));
 sky130_fd_sc_hd__nand2_1 _21609_ (.A(_05651_),
    .B(_04104_),
    .Y(_05652_));
 sky130_fd_sc_hd__a21bo_1 _21610_ (.A1(_05652_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_05653_));
 sky130_fd_sc_hd__clkbuf_8 _21611_ (.A(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__mux2_1 _21612_ (.A0(_05318_),
    .A1(net2845),
    .S(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__clkbuf_1 _21613_ (.A(_05655_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _21614_ (.A0(_05324_),
    .A1(net3325),
    .S(_05654_),
    .X(_05656_));
 sky130_fd_sc_hd__clkbuf_1 _21615_ (.A(_05656_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _21616_ (.A0(_05326_),
    .A1(net3716),
    .S(_05654_),
    .X(_05657_));
 sky130_fd_sc_hd__clkbuf_1 _21617_ (.A(_05657_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _21618_ (.A0(_05328_),
    .A1(net2635),
    .S(_05654_),
    .X(_05658_));
 sky130_fd_sc_hd__clkbuf_1 _21619_ (.A(_05658_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _21620_ (.A0(_05330_),
    .A1(net2587),
    .S(_05654_),
    .X(_05659_));
 sky130_fd_sc_hd__clkbuf_1 _21621_ (.A(_05659_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _21622_ (.A0(_05332_),
    .A1(net3374),
    .S(_05654_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _21623_ (.A(_05660_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _21624_ (.A0(_05334_),
    .A1(net3637),
    .S(_05654_),
    .X(_05661_));
 sky130_fd_sc_hd__clkbuf_1 _21625_ (.A(_05661_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _21626_ (.A0(_05336_),
    .A1(net2829),
    .S(_05654_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _21627_ (.A(_05662_),
    .X(_01338_));
 sky130_fd_sc_hd__buf_4 _21628_ (.A(_05652_),
    .X(_05663_));
 sky130_fd_sc_hd__buf_4 _21629_ (.A(_05183_),
    .X(_05664_));
 sky130_fd_sc_hd__buf_4 _21630_ (.A(_05652_),
    .X(_05665_));
 sky130_fd_sc_hd__nand2_1 _21631_ (.A(_05665_),
    .B(_05010_),
    .Y(_05666_));
 sky130_fd_sc_hd__o211a_1 _21632_ (.A1(_05095_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _21633_ (.A0(_05667_),
    .A1(net2169),
    .S(_05654_),
    .X(_05668_));
 sky130_fd_sc_hd__clkbuf_1 _21634_ (.A(_05668_),
    .X(_01339_));
 sky130_fd_sc_hd__nand2_1 _21635_ (.A(_05665_),
    .B(_05014_),
    .Y(_05669_));
 sky130_fd_sc_hd__o211a_1 _21636_ (.A1(_05101_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_1 _21637_ (.A0(_05670_),
    .A1(net2795),
    .S(_05654_),
    .X(_05671_));
 sky130_fd_sc_hd__clkbuf_1 _21638_ (.A(_05671_),
    .X(_01340_));
 sky130_fd_sc_hd__nand2_1 _21639_ (.A(_05665_),
    .B(_05018_),
    .Y(_05672_));
 sky130_fd_sc_hd__o211a_1 _21640_ (.A1(_05105_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _21641_ (.A0(_05673_),
    .A1(net3644),
    .S(_05654_),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_1 _21642_ (.A(_05674_),
    .X(_01341_));
 sky130_fd_sc_hd__nand2_1 _21643_ (.A(_05665_),
    .B(_05022_),
    .Y(_05675_));
 sky130_fd_sc_hd__o211a_1 _21644_ (.A1(_05109_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__mux2_1 _21645_ (.A0(_05676_),
    .A1(net2937),
    .S(_05654_),
    .X(_05677_));
 sky130_fd_sc_hd__clkbuf_1 _21646_ (.A(_05677_),
    .X(_01342_));
 sky130_fd_sc_hd__nand2_1 _21647_ (.A(_05665_),
    .B(_05026_),
    .Y(_05678_));
 sky130_fd_sc_hd__o211a_1 _21648_ (.A1(_05113_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _21649_ (.A0(_05679_),
    .A1(net3093),
    .S(_05654_),
    .X(_05680_));
 sky130_fd_sc_hd__clkbuf_1 _21650_ (.A(_05680_),
    .X(_01343_));
 sky130_fd_sc_hd__nand2_1 _21651_ (.A(_05665_),
    .B(_05030_),
    .Y(_05681_));
 sky130_fd_sc_hd__o211a_1 _21652_ (.A1(_05117_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _21653_ (.A0(_05682_),
    .A1(net2837),
    .S(_05654_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_1 _21654_ (.A(_05683_),
    .X(_01344_));
 sky130_fd_sc_hd__nand2_1 _21655_ (.A(_05665_),
    .B(_05034_),
    .Y(_05684_));
 sky130_fd_sc_hd__o211a_1 _21656_ (.A1(_05121_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__mux2_1 _21657_ (.A0(_05685_),
    .A1(net3646),
    .S(_05654_),
    .X(_05686_));
 sky130_fd_sc_hd__clkbuf_1 _21658_ (.A(_05686_),
    .X(_01345_));
 sky130_fd_sc_hd__nand2_1 _21659_ (.A(_05665_),
    .B(_05038_),
    .Y(_05687_));
 sky130_fd_sc_hd__o211a_1 _21660_ (.A1(_05125_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_1 _21661_ (.A0(_05688_),
    .A1(net3265),
    .S(_05654_),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _21662_ (.A(_05689_),
    .X(_01346_));
 sky130_fd_sc_hd__o211a_1 _21663_ (.A1(_05129_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05666_),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_8 _21664_ (.A(_05653_),
    .X(_05691_));
 sky130_fd_sc_hd__mux2_1 _21665_ (.A0(_05690_),
    .A1(net2704),
    .S(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__clkbuf_1 _21666_ (.A(_05692_),
    .X(_01347_));
 sky130_fd_sc_hd__o211a_1 _21667_ (.A1(_05134_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05669_),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_1 _21668_ (.A0(_05693_),
    .A1(net3151),
    .S(_05691_),
    .X(_05694_));
 sky130_fd_sc_hd__clkbuf_1 _21669_ (.A(_05694_),
    .X(_01348_));
 sky130_fd_sc_hd__o211a_1 _21670_ (.A1(_05137_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05672_),
    .X(_05695_));
 sky130_fd_sc_hd__mux2_1 _21671_ (.A0(_05695_),
    .A1(net3061),
    .S(_05691_),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_1 _21672_ (.A(_05696_),
    .X(_01349_));
 sky130_fd_sc_hd__o211a_1 _21673_ (.A1(_05140_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05675_),
    .X(_05697_));
 sky130_fd_sc_hd__mux2_1 _21674_ (.A0(_05697_),
    .A1(net3337),
    .S(_05691_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _21675_ (.A(_05698_),
    .X(_01350_));
 sky130_fd_sc_hd__o211a_1 _21676_ (.A1(_05143_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05678_),
    .X(_05699_));
 sky130_fd_sc_hd__mux2_1 _21677_ (.A0(_05699_),
    .A1(net3368),
    .S(_05691_),
    .X(_05700_));
 sky130_fd_sc_hd__clkbuf_1 _21678_ (.A(_05700_),
    .X(_01351_));
 sky130_fd_sc_hd__o211a_1 _21679_ (.A1(_05146_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05681_),
    .X(_05701_));
 sky130_fd_sc_hd__mux2_1 _21680_ (.A0(_05701_),
    .A1(net2593),
    .S(_05691_),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_1 _21681_ (.A(_05702_),
    .X(_01352_));
 sky130_fd_sc_hd__o211a_1 _21682_ (.A1(_05149_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05684_),
    .X(_05703_));
 sky130_fd_sc_hd__mux2_1 _21683_ (.A0(_05703_),
    .A1(net2930),
    .S(_05691_),
    .X(_05704_));
 sky130_fd_sc_hd__clkbuf_1 _21684_ (.A(_05704_),
    .X(_01353_));
 sky130_fd_sc_hd__o211a_1 _21685_ (.A1(_05152_),
    .A2(_05663_),
    .B1(_05664_),
    .C1(_05687_),
    .X(_05705_));
 sky130_fd_sc_hd__mux2_1 _21686_ (.A0(_05705_),
    .A1(net3101),
    .S(_05691_),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_1 _21687_ (.A(_05706_),
    .X(_01354_));
 sky130_fd_sc_hd__clkbuf_8 _21688_ (.A(_05183_),
    .X(_05707_));
 sky130_fd_sc_hd__o211a_1 _21689_ (.A1(_05059_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05666_),
    .X(_05708_));
 sky130_fd_sc_hd__mux2_1 _21690_ (.A0(_05708_),
    .A1(net2346),
    .S(_05691_),
    .X(_05709_));
 sky130_fd_sc_hd__clkbuf_1 _21691_ (.A(_05709_),
    .X(_01355_));
 sky130_fd_sc_hd__o211a_1 _21692_ (.A1(_05063_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05669_),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_1 _21693_ (.A0(_05710_),
    .A1(net3566),
    .S(_05691_),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _21694_ (.A(_05711_),
    .X(_01356_));
 sky130_fd_sc_hd__o211a_1 _21695_ (.A1(_05066_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05672_),
    .X(_05712_));
 sky130_fd_sc_hd__mux2_1 _21696_ (.A0(_05712_),
    .A1(net2410),
    .S(_05691_),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_1 _21697_ (.A(_05713_),
    .X(_01357_));
 sky130_fd_sc_hd__o211a_1 _21698_ (.A1(_05069_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05675_),
    .X(_05714_));
 sky130_fd_sc_hd__mux2_1 _21699_ (.A0(_05714_),
    .A1(net2792),
    .S(_05691_),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_1 _21700_ (.A(_05715_),
    .X(_01358_));
 sky130_fd_sc_hd__o211a_1 _21701_ (.A1(_05072_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05678_),
    .X(_05716_));
 sky130_fd_sc_hd__mux2_1 _21702_ (.A0(_05716_),
    .A1(net2366),
    .S(_05691_),
    .X(_05717_));
 sky130_fd_sc_hd__clkbuf_1 _21703_ (.A(_05717_),
    .X(_01359_));
 sky130_fd_sc_hd__o211a_1 _21704_ (.A1(_05075_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05681_),
    .X(_05718_));
 sky130_fd_sc_hd__mux2_1 _21705_ (.A0(_05718_),
    .A1(net3398),
    .S(_05691_),
    .X(_05719_));
 sky130_fd_sc_hd__clkbuf_1 _21706_ (.A(_05719_),
    .X(_01360_));
 sky130_fd_sc_hd__o211a_1 _21707_ (.A1(_05078_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05684_),
    .X(_05720_));
 sky130_fd_sc_hd__mux2_1 _21708_ (.A0(_05720_),
    .A1(net2895),
    .S(_05691_),
    .X(_05721_));
 sky130_fd_sc_hd__clkbuf_1 _21709_ (.A(_05721_),
    .X(_01361_));
 sky130_fd_sc_hd__o211a_1 _21710_ (.A1(_05081_),
    .A2(_05665_),
    .B1(_05707_),
    .C1(_05687_),
    .X(_05722_));
 sky130_fd_sc_hd__mux2_1 _21711_ (.A0(_05722_),
    .A1(net2788),
    .S(_05691_),
    .X(_05723_));
 sky130_fd_sc_hd__clkbuf_1 _21712_ (.A(_05723_),
    .X(_01362_));
 sky130_fd_sc_hd__nand2_1 _21713_ (.A(_05651_),
    .B(_04183_),
    .Y(_05724_));
 sky130_fd_sc_hd__inv_2 _21714_ (.A(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_4 _21715_ (.A1(_05471_),
    .A2(_05725_),
    .B1(_04776_),
    .Y(_05726_));
 sky130_fd_sc_hd__mux2_1 _21716_ (.A0(_05318_),
    .A1(net3706),
    .S(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _21717_ (.A(_05727_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _21718_ (.A0(_05324_),
    .A1(net2420),
    .S(_05726_),
    .X(_05728_));
 sky130_fd_sc_hd__clkbuf_1 _21719_ (.A(_05728_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _21720_ (.A0(_05326_),
    .A1(net3593),
    .S(_05726_),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _21721_ (.A(_05729_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _21722_ (.A0(_05328_),
    .A1(net2273),
    .S(_05726_),
    .X(_05730_));
 sky130_fd_sc_hd__clkbuf_1 _21723_ (.A(_05730_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _21724_ (.A0(_05330_),
    .A1(net2217),
    .S(_05726_),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_1 _21725_ (.A(_05731_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _21726_ (.A0(_05332_),
    .A1(net2431),
    .S(_05726_),
    .X(_05732_));
 sky130_fd_sc_hd__clkbuf_1 _21727_ (.A(_05732_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _21728_ (.A0(_05334_),
    .A1(net2826),
    .S(_05726_),
    .X(_05733_));
 sky130_fd_sc_hd__clkbuf_1 _21729_ (.A(_05733_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _21730_ (.A0(_05336_),
    .A1(net2463),
    .S(_05726_),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_1 _21731_ (.A(_05734_),
    .X(_01370_));
 sky130_fd_sc_hd__buf_4 _21732_ (.A(_05726_),
    .X(_05735_));
 sky130_fd_sc_hd__buf_4 _21733_ (.A(_05725_),
    .X(_05736_));
 sky130_fd_sc_hd__buf_4 _21734_ (.A(_05725_),
    .X(_05737_));
 sky130_fd_sc_hd__nor2_1 _21735_ (.A(_05583_),
    .B(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__a211o_1 _21736_ (.A1(_05484_),
    .A2(_05736_),
    .B1(_05622_),
    .C1(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__buf_4 _21737_ (.A(_05726_),
    .X(_05740_));
 sky130_fd_sc_hd__nand2_1 _21738_ (.A(_05740_),
    .B(net1951),
    .Y(_05741_));
 sky130_fd_sc_hd__o21ai_1 _21739_ (.A1(_05735_),
    .A2(_05739_),
    .B1(_05741_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _21740_ (.A(_05589_),
    .B(_05737_),
    .Y(_05742_));
 sky130_fd_sc_hd__a211o_1 _21741_ (.A1(_05491_),
    .A2(_05736_),
    .B1(_05622_),
    .C1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__nand2_1 _21742_ (.A(_05740_),
    .B(net1466),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_1 _21743_ (.A1(_05735_),
    .A2(_05743_),
    .B1(net1467),
    .Y(_01372_));
 sky130_fd_sc_hd__buf_4 _21744_ (.A(_04598_),
    .X(_05745_));
 sky130_fd_sc_hd__nor2_1 _21745_ (.A(_05593_),
    .B(_05737_),
    .Y(_05746_));
 sky130_fd_sc_hd__a211o_1 _21746_ (.A1(_05495_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__nand2_1 _21747_ (.A(_05740_),
    .B(net1958),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_1 _21748_ (.A1(_05735_),
    .A2(_05747_),
    .B1(_05748_),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_1 _21749_ (.A(_05597_),
    .B(_05737_),
    .Y(_05749_));
 sky130_fd_sc_hd__a211o_1 _21750_ (.A1(_05500_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__nand2_1 _21751_ (.A(_05740_),
    .B(net1508),
    .Y(_05751_));
 sky130_fd_sc_hd__o21ai_1 _21752_ (.A1(_05735_),
    .A2(_05750_),
    .B1(net1509),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _21753_ (.A(_05601_),
    .B(_05737_),
    .Y(_05752_));
 sky130_fd_sc_hd__a211o_1 _21754_ (.A1(_05504_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2_1 _21755_ (.A(_05740_),
    .B(net1554),
    .Y(_05754_));
 sky130_fd_sc_hd__o21ai_1 _21756_ (.A1(_05735_),
    .A2(_05753_),
    .B1(net1555),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_1 _21757_ (.A(_05605_),
    .B(_05737_),
    .Y(_05755_));
 sky130_fd_sc_hd__a211o_1 _21758_ (.A1(_05508_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__nand2_1 _21759_ (.A(_05740_),
    .B(net1832),
    .Y(_05757_));
 sky130_fd_sc_hd__o21ai_1 _21760_ (.A1(_05735_),
    .A2(_05756_),
    .B1(net1833),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _21761_ (.A(_05609_),
    .B(_05737_),
    .Y(_05758_));
 sky130_fd_sc_hd__a211o_1 _21762_ (.A1(_05512_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__nand2_1 _21763_ (.A(_05740_),
    .B(net1080),
    .Y(_05760_));
 sky130_fd_sc_hd__o21ai_1 _21764_ (.A1(_05735_),
    .A2(_05759_),
    .B1(net1081),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _21765_ (.A(_05613_),
    .B(_05737_),
    .Y(_05761_));
 sky130_fd_sc_hd__a211o_1 _21766_ (.A1(_05516_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__nand2_1 _21767_ (.A(_05740_),
    .B(net832),
    .Y(_05763_));
 sky130_fd_sc_hd__o21ai_1 _21768_ (.A1(_05735_),
    .A2(_05762_),
    .B1(net833),
    .Y(_01378_));
 sky130_fd_sc_hd__buf_4 _21769_ (.A(_05726_),
    .X(_05764_));
 sky130_fd_sc_hd__a211o_1 _21770_ (.A1(_05521_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05738_),
    .X(_05765_));
 sky130_fd_sc_hd__nand2_1 _21771_ (.A(_05740_),
    .B(net844),
    .Y(_05766_));
 sky130_fd_sc_hd__o21ai_1 _21772_ (.A1(_05764_),
    .A2(_05765_),
    .B1(net845),
    .Y(_01379_));
 sky130_fd_sc_hd__a211o_1 _21773_ (.A1(_05524_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05742_),
    .X(_05767_));
 sky130_fd_sc_hd__nand2_1 _21774_ (.A(_05740_),
    .B(net1270),
    .Y(_05768_));
 sky130_fd_sc_hd__o21ai_1 _21775_ (.A1(_05764_),
    .A2(_05767_),
    .B1(net1271),
    .Y(_01380_));
 sky130_fd_sc_hd__a211o_1 _21776_ (.A1(_05527_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05746_),
    .X(_05769_));
 sky130_fd_sc_hd__nand2_1 _21777_ (.A(_05740_),
    .B(net900),
    .Y(_05770_));
 sky130_fd_sc_hd__o21ai_1 _21778_ (.A1(_05764_),
    .A2(_05769_),
    .B1(net901),
    .Y(_01381_));
 sky130_fd_sc_hd__a211o_1 _21779_ (.A1(_05530_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05749_),
    .X(_05771_));
 sky130_fd_sc_hd__nand2_1 _21780_ (.A(_05740_),
    .B(net1768),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_1 _21781_ (.A1(_05764_),
    .A2(_05771_),
    .B1(net1769),
    .Y(_01382_));
 sky130_fd_sc_hd__a211o_1 _21782_ (.A1(_05533_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05752_),
    .X(_05773_));
 sky130_fd_sc_hd__nand2_1 _21783_ (.A(_05740_),
    .B(net1410),
    .Y(_05774_));
 sky130_fd_sc_hd__o21ai_1 _21784_ (.A1(_05764_),
    .A2(_05773_),
    .B1(net1411),
    .Y(_01383_));
 sky130_fd_sc_hd__a211o_1 _21785_ (.A1(_05536_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05755_),
    .X(_05775_));
 sky130_fd_sc_hd__nand2_1 _21786_ (.A(_05740_),
    .B(net1478),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_1 _21787_ (.A1(_05764_),
    .A2(_05775_),
    .B1(net1479),
    .Y(_01384_));
 sky130_fd_sc_hd__a211o_1 _21788_ (.A1(_05539_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05758_),
    .X(_05777_));
 sky130_fd_sc_hd__nand2_1 _21789_ (.A(_05740_),
    .B(net802),
    .Y(_05778_));
 sky130_fd_sc_hd__o21ai_1 _21790_ (.A1(_05764_),
    .A2(_05777_),
    .B1(net803),
    .Y(_01385_));
 sky130_fd_sc_hd__a211o_1 _21791_ (.A1(_05542_),
    .A2(_05736_),
    .B1(_05745_),
    .C1(_05761_),
    .X(_05779_));
 sky130_fd_sc_hd__nand2_1 _21792_ (.A(_05740_),
    .B(net868),
    .Y(_05780_));
 sky130_fd_sc_hd__o21ai_1 _21793_ (.A1(_05764_),
    .A2(_05779_),
    .B1(net869),
    .Y(_01386_));
 sky130_fd_sc_hd__a211o_1 _21794_ (.A1(_05545_),
    .A2(_05737_),
    .B1(_05745_),
    .C1(_05738_),
    .X(_05781_));
 sky130_fd_sc_hd__nand2_1 _21795_ (.A(_05735_),
    .B(net1088),
    .Y(_05782_));
 sky130_fd_sc_hd__o21ai_1 _21796_ (.A1(_05764_),
    .A2(_05781_),
    .B1(net1089),
    .Y(_01387_));
 sky130_fd_sc_hd__a211o_1 _21797_ (.A1(_05548_),
    .A2(_05737_),
    .B1(_05745_),
    .C1(_05742_),
    .X(_05783_));
 sky130_fd_sc_hd__nand2_1 _21798_ (.A(_05735_),
    .B(net1248),
    .Y(_05784_));
 sky130_fd_sc_hd__o21ai_1 _21799_ (.A1(_05764_),
    .A2(_05783_),
    .B1(net1249),
    .Y(_01388_));
 sky130_fd_sc_hd__buf_4 _21800_ (.A(_04598_),
    .X(_05785_));
 sky130_fd_sc_hd__a211o_1 _21801_ (.A1(_05551_),
    .A2(_05737_),
    .B1(_05785_),
    .C1(_05746_),
    .X(_05786_));
 sky130_fd_sc_hd__nand2_1 _21802_ (.A(_05735_),
    .B(net1646),
    .Y(_05787_));
 sky130_fd_sc_hd__o21ai_1 _21803_ (.A1(_05764_),
    .A2(_05786_),
    .B1(net1647),
    .Y(_01389_));
 sky130_fd_sc_hd__a211o_1 _21804_ (.A1(_05555_),
    .A2(_05737_),
    .B1(_05785_),
    .C1(_05749_),
    .X(_05788_));
 sky130_fd_sc_hd__nand2_1 _21805_ (.A(_05735_),
    .B(net1092),
    .Y(_05789_));
 sky130_fd_sc_hd__o21ai_1 _21806_ (.A1(_05764_),
    .A2(_05788_),
    .B1(net1093),
    .Y(_01390_));
 sky130_fd_sc_hd__a211o_1 _21807_ (.A1(_05558_),
    .A2(_05737_),
    .B1(_05785_),
    .C1(_05752_),
    .X(_05790_));
 sky130_fd_sc_hd__nand2_1 _21808_ (.A(_05735_),
    .B(net1424),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_1 _21809_ (.A1(_05764_),
    .A2(_05790_),
    .B1(net1425),
    .Y(_01391_));
 sky130_fd_sc_hd__a211o_1 _21810_ (.A1(_05561_),
    .A2(_05737_),
    .B1(_05785_),
    .C1(_05755_),
    .X(_05792_));
 sky130_fd_sc_hd__nand2_1 _21811_ (.A(_05735_),
    .B(net1074),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_1 _21812_ (.A1(_05764_),
    .A2(_05792_),
    .B1(net1075),
    .Y(_01392_));
 sky130_fd_sc_hd__a211o_1 _21813_ (.A1(_05564_),
    .A2(_05737_),
    .B1(_05785_),
    .C1(_05758_),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_1 _21814_ (.A(_05735_),
    .B(net1064),
    .Y(_05795_));
 sky130_fd_sc_hd__o21ai_1 _21815_ (.A1(_05764_),
    .A2(_05794_),
    .B1(net1065),
    .Y(_01393_));
 sky130_fd_sc_hd__a211o_1 _21816_ (.A1(_05567_),
    .A2(_05737_),
    .B1(_05785_),
    .C1(_05761_),
    .X(_05796_));
 sky130_fd_sc_hd__nand2_1 _21817_ (.A(_05735_),
    .B(net1718),
    .Y(_05797_));
 sky130_fd_sc_hd__o21ai_1 _21818_ (.A1(_05764_),
    .A2(_05796_),
    .B1(net1719),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_1 _21819_ (.A(_05651_),
    .B(_04257_),
    .Y(_05798_));
 sky130_fd_sc_hd__inv_2 _21820_ (.A(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_4 _21821_ (.A1(_05471_),
    .A2(_05799_),
    .B1(_04776_),
    .Y(_05800_));
 sky130_fd_sc_hd__mux2_1 _21822_ (.A0(_05318_),
    .A1(net3615),
    .S(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_1 _21823_ (.A(_05801_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _21824_ (.A0(_05324_),
    .A1(net2617),
    .S(_05800_),
    .X(_05802_));
 sky130_fd_sc_hd__clkbuf_1 _21825_ (.A(_05802_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _21826_ (.A0(_05326_),
    .A1(net3718),
    .S(_05800_),
    .X(_05803_));
 sky130_fd_sc_hd__clkbuf_1 _21827_ (.A(_05803_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _21828_ (.A0(_05328_),
    .A1(net3306),
    .S(_05800_),
    .X(_05804_));
 sky130_fd_sc_hd__clkbuf_1 _21829_ (.A(_05804_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _21830_ (.A0(_05330_),
    .A1(net2639),
    .S(_05800_),
    .X(_05805_));
 sky130_fd_sc_hd__clkbuf_1 _21831_ (.A(_05805_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _21832_ (.A0(_05332_),
    .A1(net2206),
    .S(_05800_),
    .X(_05806_));
 sky130_fd_sc_hd__clkbuf_1 _21833_ (.A(_05806_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _21834_ (.A0(_05334_),
    .A1(net2369),
    .S(_05800_),
    .X(_05807_));
 sky130_fd_sc_hd__clkbuf_1 _21835_ (.A(_05807_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _21836_ (.A0(_05336_),
    .A1(net2715),
    .S(_05800_),
    .X(_05808_));
 sky130_fd_sc_hd__clkbuf_1 _21837_ (.A(_05808_),
    .X(_01402_));
 sky130_fd_sc_hd__buf_4 _21838_ (.A(_05800_),
    .X(_05809_));
 sky130_fd_sc_hd__buf_4 _21839_ (.A(_05799_),
    .X(_05810_));
 sky130_fd_sc_hd__buf_4 _21840_ (.A(_05799_),
    .X(_05811_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(_05583_),
    .B(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__a211o_1 _21842_ (.A1(_05484_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__buf_4 _21843_ (.A(_05800_),
    .X(_05814_));
 sky130_fd_sc_hd__nand2_1 _21844_ (.A(_05814_),
    .B(net1967),
    .Y(_05815_));
 sky130_fd_sc_hd__o21ai_1 _21845_ (.A1(_05809_),
    .A2(_05813_),
    .B1(_05815_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor2_1 _21846_ (.A(_05589_),
    .B(_05811_),
    .Y(_05816_));
 sky130_fd_sc_hd__a211o_1 _21847_ (.A1(_05491_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_1 _21848_ (.A(_05814_),
    .B(net1704),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_1 _21849_ (.A1(_05809_),
    .A2(_05817_),
    .B1(net1705),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_1 _21850_ (.A(_05593_),
    .B(_05811_),
    .Y(_05819_));
 sky130_fd_sc_hd__a211o_1 _21851_ (.A1(_05495_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__nand2_1 _21852_ (.A(_05814_),
    .B(net1893),
    .Y(_05821_));
 sky130_fd_sc_hd__o21ai_1 _21853_ (.A1(_05809_),
    .A2(_05820_),
    .B1(net1894),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _21854_ (.A(_05597_),
    .B(_05811_),
    .Y(_05822_));
 sky130_fd_sc_hd__a211o_1 _21855_ (.A1(_05500_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__nand2_1 _21856_ (.A(_05814_),
    .B(net940),
    .Y(_05824_));
 sky130_fd_sc_hd__o21ai_1 _21857_ (.A1(_05809_),
    .A2(_05823_),
    .B1(net941),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _21858_ (.A(_05601_),
    .B(_05811_),
    .Y(_05825_));
 sky130_fd_sc_hd__a211o_1 _21859_ (.A1(_05504_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05825_),
    .X(_05826_));
 sky130_fd_sc_hd__nand2_1 _21860_ (.A(_05814_),
    .B(net1638),
    .Y(_05827_));
 sky130_fd_sc_hd__o21ai_1 _21861_ (.A1(_05809_),
    .A2(_05826_),
    .B1(net1639),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(_05605_),
    .B(_05811_),
    .Y(_05828_));
 sky130_fd_sc_hd__a211o_1 _21863_ (.A1(_05508_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__nand2_1 _21864_ (.A(_05814_),
    .B(net1562),
    .Y(_05830_));
 sky130_fd_sc_hd__o21ai_1 _21865_ (.A1(_05809_),
    .A2(_05829_),
    .B1(net1563),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_1 _21866_ (.A(_05609_),
    .B(_05811_),
    .Y(_05831_));
 sky130_fd_sc_hd__a211o_1 _21867_ (.A1(_05512_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__nand2_1 _21868_ (.A(_05814_),
    .B(net1200),
    .Y(_05833_));
 sky130_fd_sc_hd__o21ai_1 _21869_ (.A1(_05809_),
    .A2(_05832_),
    .B1(net1201),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _21870_ (.A(_05613_),
    .B(_05811_),
    .Y(_05834_));
 sky130_fd_sc_hd__a211o_1 _21871_ (.A1(_05516_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__nand2_1 _21872_ (.A(_05814_),
    .B(net1392),
    .Y(_05836_));
 sky130_fd_sc_hd__o21ai_1 _21873_ (.A1(_05809_),
    .A2(_05835_),
    .B1(net1393),
    .Y(_01410_));
 sky130_fd_sc_hd__buf_4 _21874_ (.A(_05800_),
    .X(_05837_));
 sky130_fd_sc_hd__a211o_1 _21875_ (.A1(_05521_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05812_),
    .X(_05838_));
 sky130_fd_sc_hd__nand2_1 _21876_ (.A(_05814_),
    .B(net1879),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_1 _21877_ (.A1(_05837_),
    .A2(_05838_),
    .B1(net1880),
    .Y(_01411_));
 sky130_fd_sc_hd__a211o_1 _21878_ (.A1(_05524_),
    .A2(_05810_),
    .B1(_05785_),
    .C1(_05816_),
    .X(_05840_));
 sky130_fd_sc_hd__nand2_1 _21879_ (.A(_05814_),
    .B(net1826),
    .Y(_05841_));
 sky130_fd_sc_hd__o21ai_1 _21880_ (.A1(_05837_),
    .A2(_05840_),
    .B1(net1827),
    .Y(_01412_));
 sky130_fd_sc_hd__buf_4 _21881_ (.A(_04598_),
    .X(_05842_));
 sky130_fd_sc_hd__a211o_1 _21882_ (.A1(_05527_),
    .A2(_05810_),
    .B1(_05842_),
    .C1(_05819_),
    .X(_05843_));
 sky130_fd_sc_hd__nand2_1 _21883_ (.A(_05814_),
    .B(net1686),
    .Y(_05844_));
 sky130_fd_sc_hd__o21ai_1 _21884_ (.A1(_05837_),
    .A2(_05843_),
    .B1(net1687),
    .Y(_01413_));
 sky130_fd_sc_hd__a211o_1 _21885_ (.A1(_05530_),
    .A2(_05810_),
    .B1(_05842_),
    .C1(_05822_),
    .X(_05845_));
 sky130_fd_sc_hd__nand2_1 _21886_ (.A(_05814_),
    .B(net974),
    .Y(_05846_));
 sky130_fd_sc_hd__o21ai_1 _21887_ (.A1(_05837_),
    .A2(_05845_),
    .B1(net975),
    .Y(_01414_));
 sky130_fd_sc_hd__a211o_1 _21888_ (.A1(_05533_),
    .A2(_05810_),
    .B1(_05842_),
    .C1(_05825_),
    .X(_05847_));
 sky130_fd_sc_hd__nand2_1 _21889_ (.A(_05814_),
    .B(net1104),
    .Y(_05848_));
 sky130_fd_sc_hd__o21ai_1 _21890_ (.A1(_05837_),
    .A2(_05847_),
    .B1(net1105),
    .Y(_01415_));
 sky130_fd_sc_hd__a211o_1 _21891_ (.A1(_05536_),
    .A2(_05810_),
    .B1(_05842_),
    .C1(_05828_),
    .X(_05849_));
 sky130_fd_sc_hd__nand2_1 _21892_ (.A(_05814_),
    .B(net1440),
    .Y(_05850_));
 sky130_fd_sc_hd__o21ai_1 _21893_ (.A1(_05837_),
    .A2(_05849_),
    .B1(net1441),
    .Y(_01416_));
 sky130_fd_sc_hd__a211o_1 _21894_ (.A1(_05539_),
    .A2(_05810_),
    .B1(_05842_),
    .C1(_05831_),
    .X(_05851_));
 sky130_fd_sc_hd__nand2_1 _21895_ (.A(_05814_),
    .B(net1364),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ai_1 _21896_ (.A1(_05837_),
    .A2(_05851_),
    .B1(net1365),
    .Y(_01417_));
 sky130_fd_sc_hd__a211o_1 _21897_ (.A1(_05542_),
    .A2(_05810_),
    .B1(_05842_),
    .C1(_05834_),
    .X(_05853_));
 sky130_fd_sc_hd__nand2_1 _21898_ (.A(_05814_),
    .B(net1909),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_1 _21899_ (.A1(_05837_),
    .A2(_05853_),
    .B1(net1910),
    .Y(_01418_));
 sky130_fd_sc_hd__a211o_1 _21900_ (.A1(_05545_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05812_),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _21901_ (.A(_05809_),
    .B(net708),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_1 _21902_ (.A1(_05837_),
    .A2(_05855_),
    .B1(net709),
    .Y(_01419_));
 sky130_fd_sc_hd__a211o_1 _21903_ (.A1(_05548_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05816_),
    .X(_05857_));
 sky130_fd_sc_hd__nand2_1 _21904_ (.A(_05809_),
    .B(net1318),
    .Y(_05858_));
 sky130_fd_sc_hd__o21ai_1 _21905_ (.A1(_05837_),
    .A2(_05857_),
    .B1(net1319),
    .Y(_01420_));
 sky130_fd_sc_hd__a211o_1 _21906_ (.A1(_05551_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05819_),
    .X(_05859_));
 sky130_fd_sc_hd__nand2_1 _21907_ (.A(_05809_),
    .B(net744),
    .Y(_05860_));
 sky130_fd_sc_hd__o21ai_1 _21908_ (.A1(_05837_),
    .A2(_05859_),
    .B1(net745),
    .Y(_01421_));
 sky130_fd_sc_hd__a211o_1 _21909_ (.A1(_05555_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05822_),
    .X(_05861_));
 sky130_fd_sc_hd__nand2_1 _21910_ (.A(_05809_),
    .B(net1224),
    .Y(_05862_));
 sky130_fd_sc_hd__o21ai_1 _21911_ (.A1(_05837_),
    .A2(_05861_),
    .B1(net1225),
    .Y(_01422_));
 sky130_fd_sc_hd__a211o_1 _21912_ (.A1(_05558_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05825_),
    .X(_05863_));
 sky130_fd_sc_hd__nand2_1 _21913_ (.A(_05809_),
    .B(net1504),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_1 _21914_ (.A1(_05837_),
    .A2(_05863_),
    .B1(net1505),
    .Y(_01423_));
 sky130_fd_sc_hd__a211o_1 _21915_ (.A1(_05561_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05828_),
    .X(_05865_));
 sky130_fd_sc_hd__nand2_1 _21916_ (.A(_05809_),
    .B(net1484),
    .Y(_05866_));
 sky130_fd_sc_hd__o21ai_1 _21917_ (.A1(_05837_),
    .A2(_05865_),
    .B1(net1485),
    .Y(_01424_));
 sky130_fd_sc_hd__a211o_1 _21918_ (.A1(_05564_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05831_),
    .X(_05867_));
 sky130_fd_sc_hd__nand2_1 _21919_ (.A(_05809_),
    .B(net1246),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_1 _21920_ (.A1(_05837_),
    .A2(_05867_),
    .B1(net1247),
    .Y(_01425_));
 sky130_fd_sc_hd__a211o_1 _21921_ (.A1(_05567_),
    .A2(_05811_),
    .B1(_05842_),
    .C1(_05834_),
    .X(_05869_));
 sky130_fd_sc_hd__nand2_1 _21922_ (.A(_05809_),
    .B(net1782),
    .Y(_05870_));
 sky130_fd_sc_hd__o21ai_1 _21923_ (.A1(_05837_),
    .A2(_05869_),
    .B1(net1783),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _21924_ (.A(_05651_),
    .B(_04333_),
    .Y(_05871_));
 sky130_fd_sc_hd__inv_2 _21925_ (.A(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_4 _21926_ (.A1(_05471_),
    .A2(_05872_),
    .B1(_04776_),
    .Y(_05873_));
 sky130_fd_sc_hd__mux2_1 _21927_ (.A0(_05318_),
    .A1(net2675),
    .S(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__clkbuf_1 _21928_ (.A(_05874_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _21929_ (.A0(_05324_),
    .A1(net2972),
    .S(_05873_),
    .X(_05875_));
 sky130_fd_sc_hd__clkbuf_1 _21930_ (.A(_05875_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _21931_ (.A0(_05326_),
    .A1(net2847),
    .S(_05873_),
    .X(_05876_));
 sky130_fd_sc_hd__clkbuf_1 _21932_ (.A(_05876_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _21933_ (.A0(_05328_),
    .A1(net3327),
    .S(_05873_),
    .X(_05877_));
 sky130_fd_sc_hd__clkbuf_1 _21934_ (.A(_05877_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _21935_ (.A0(_05330_),
    .A1(net2201),
    .S(_05873_),
    .X(_05878_));
 sky130_fd_sc_hd__clkbuf_1 _21936_ (.A(_05878_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _21937_ (.A0(_05332_),
    .A1(net3597),
    .S(_05873_),
    .X(_05879_));
 sky130_fd_sc_hd__clkbuf_1 _21938_ (.A(_05879_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _21939_ (.A0(_05334_),
    .A1(net2804),
    .S(_05873_),
    .X(_05880_));
 sky130_fd_sc_hd__clkbuf_1 _21940_ (.A(_05880_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _21941_ (.A0(_05336_),
    .A1(net3677),
    .S(_05873_),
    .X(_05881_));
 sky130_fd_sc_hd__clkbuf_1 _21942_ (.A(_05881_),
    .X(_01434_));
 sky130_fd_sc_hd__buf_4 _21943_ (.A(_05873_),
    .X(_05882_));
 sky130_fd_sc_hd__buf_4 _21944_ (.A(_05872_),
    .X(_05883_));
 sky130_fd_sc_hd__buf_4 _21945_ (.A(_05872_),
    .X(_05884_));
 sky130_fd_sc_hd__nor2_1 _21946_ (.A(_05583_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__a211o_1 _21947_ (.A1(_05484_),
    .A2(_05883_),
    .B1(_05842_),
    .C1(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__buf_4 _21948_ (.A(_05873_),
    .X(_05887_));
 sky130_fd_sc_hd__nand2_1 _21949_ (.A(_05887_),
    .B(net1192),
    .Y(_05888_));
 sky130_fd_sc_hd__o21ai_1 _21950_ (.A1(_05882_),
    .A2(_05886_),
    .B1(net1193),
    .Y(_01435_));
 sky130_fd_sc_hd__nor2_1 _21951_ (.A(_05589_),
    .B(_05884_),
    .Y(_05889_));
 sky130_fd_sc_hd__a211o_1 _21952_ (.A1(_05491_),
    .A2(_05883_),
    .B1(_05842_),
    .C1(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__nand2_1 _21953_ (.A(_05887_),
    .B(net1368),
    .Y(_05891_));
 sky130_fd_sc_hd__o21ai_1 _21954_ (.A1(_05882_),
    .A2(_05890_),
    .B1(net1369),
    .Y(_01436_));
 sky130_fd_sc_hd__buf_8 _21955_ (.A(_09057_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_4 _21956_ (.A(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__nor2_1 _21957_ (.A(_05593_),
    .B(_05884_),
    .Y(_05894_));
 sky130_fd_sc_hd__a211o_1 _21958_ (.A1(_05495_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05894_),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_1 _21959_ (.A(_05887_),
    .B(net1030),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_1 _21960_ (.A1(_05882_),
    .A2(_05895_),
    .B1(net1031),
    .Y(_01437_));
 sky130_fd_sc_hd__nor2_1 _21961_ (.A(_05597_),
    .B(_05884_),
    .Y(_05897_));
 sky130_fd_sc_hd__a211o_1 _21962_ (.A1(_05500_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__nand2_1 _21963_ (.A(_05887_),
    .B(net892),
    .Y(_05899_));
 sky130_fd_sc_hd__o21ai_1 _21964_ (.A1(_05882_),
    .A2(_05898_),
    .B1(net893),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _21965_ (.A(_05601_),
    .B(_05884_),
    .Y(_05900_));
 sky130_fd_sc_hd__a211o_1 _21966_ (.A1(_05504_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__nand2_1 _21967_ (.A(_05887_),
    .B(net1925),
    .Y(_05902_));
 sky130_fd_sc_hd__o21ai_1 _21968_ (.A1(_05882_),
    .A2(_05901_),
    .B1(net1926),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _21969_ (.A(_05605_),
    .B(_05884_),
    .Y(_05903_));
 sky130_fd_sc_hd__a211o_1 _21970_ (.A1(_05508_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__nand2_1 _21971_ (.A(_05887_),
    .B(net796),
    .Y(_05905_));
 sky130_fd_sc_hd__o21ai_1 _21972_ (.A1(_05882_),
    .A2(_05904_),
    .B1(net797),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _21973_ (.A(_05609_),
    .B(_05884_),
    .Y(_05906_));
 sky130_fd_sc_hd__a211o_1 _21974_ (.A1(_05512_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__nand2_1 _21975_ (.A(_05887_),
    .B(net1032),
    .Y(_05908_));
 sky130_fd_sc_hd__o21ai_1 _21976_ (.A1(_05882_),
    .A2(_05907_),
    .B1(net1033),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _21977_ (.A(_05613_),
    .B(_05884_),
    .Y(_05909_));
 sky130_fd_sc_hd__a211o_1 _21978_ (.A1(_05516_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__nand2_1 _21979_ (.A(_05887_),
    .B(net1360),
    .Y(_05911_));
 sky130_fd_sc_hd__o21ai_1 _21980_ (.A1(_05882_),
    .A2(_05910_),
    .B1(net1361),
    .Y(_01442_));
 sky130_fd_sc_hd__buf_4 _21981_ (.A(_05873_),
    .X(_05912_));
 sky130_fd_sc_hd__a211o_1 _21982_ (.A1(_05521_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05885_),
    .X(_05913_));
 sky130_fd_sc_hd__nand2_1 _21983_ (.A(_05887_),
    .B(net1000),
    .Y(_05914_));
 sky130_fd_sc_hd__o21ai_1 _21984_ (.A1(_05912_),
    .A2(_05913_),
    .B1(net1001),
    .Y(_01443_));
 sky130_fd_sc_hd__a211o_1 _21985_ (.A1(_05524_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05889_),
    .X(_05915_));
 sky130_fd_sc_hd__nand2_1 _21986_ (.A(_05887_),
    .B(net1176),
    .Y(_05916_));
 sky130_fd_sc_hd__o21ai_1 _21987_ (.A1(_05912_),
    .A2(_05915_),
    .B1(net1177),
    .Y(_01444_));
 sky130_fd_sc_hd__a211o_1 _21988_ (.A1(_05527_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05894_),
    .X(_05917_));
 sky130_fd_sc_hd__nand2_1 _21989_ (.A(_05887_),
    .B(net688),
    .Y(_05918_));
 sky130_fd_sc_hd__o21ai_1 _21990_ (.A1(_05912_),
    .A2(_05917_),
    .B1(net689),
    .Y(_01445_));
 sky130_fd_sc_hd__a211o_1 _21991_ (.A1(_05530_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05897_),
    .X(_05919_));
 sky130_fd_sc_hd__nand2_1 _21992_ (.A(_05887_),
    .B(net914),
    .Y(_05920_));
 sky130_fd_sc_hd__o21ai_1 _21993_ (.A1(_05912_),
    .A2(_05919_),
    .B1(net915),
    .Y(_01446_));
 sky130_fd_sc_hd__a211o_1 _21994_ (.A1(_05533_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05900_),
    .X(_05921_));
 sky130_fd_sc_hd__nand2_1 _21995_ (.A(_05887_),
    .B(net1953),
    .Y(_05922_));
 sky130_fd_sc_hd__o21ai_1 _21996_ (.A1(_05912_),
    .A2(_05921_),
    .B1(_05922_),
    .Y(_01447_));
 sky130_fd_sc_hd__a211o_1 _21997_ (.A1(_05536_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05903_),
    .X(_05923_));
 sky130_fd_sc_hd__nand2_1 _21998_ (.A(_05887_),
    .B(net702),
    .Y(_05924_));
 sky130_fd_sc_hd__o21ai_1 _21999_ (.A1(_05912_),
    .A2(_05923_),
    .B1(net703),
    .Y(_01448_));
 sky130_fd_sc_hd__a211o_1 _22000_ (.A1(_05539_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05906_),
    .X(_05925_));
 sky130_fd_sc_hd__nand2_1 _22001_ (.A(_05887_),
    .B(net1138),
    .Y(_05926_));
 sky130_fd_sc_hd__o21ai_1 _22002_ (.A1(_05912_),
    .A2(_05925_),
    .B1(net1139),
    .Y(_01449_));
 sky130_fd_sc_hd__a211o_1 _22003_ (.A1(_05542_),
    .A2(_05883_),
    .B1(_05893_),
    .C1(_05909_),
    .X(_05927_));
 sky130_fd_sc_hd__nand2_1 _22004_ (.A(_05887_),
    .B(net1901),
    .Y(_05928_));
 sky130_fd_sc_hd__o21ai_1 _22005_ (.A1(_05912_),
    .A2(_05927_),
    .B1(net1902),
    .Y(_01450_));
 sky130_fd_sc_hd__a211o_1 _22006_ (.A1(_05545_),
    .A2(_05884_),
    .B1(_05893_),
    .C1(_05885_),
    .X(_05929_));
 sky130_fd_sc_hd__nand2_1 _22007_ (.A(_05882_),
    .B(net656),
    .Y(_05930_));
 sky130_fd_sc_hd__o21ai_1 _22008_ (.A1(_05912_),
    .A2(_05929_),
    .B1(net657),
    .Y(_01451_));
 sky130_fd_sc_hd__a211o_1 _22009_ (.A1(_05548_),
    .A2(_05884_),
    .B1(_05893_),
    .C1(_05889_),
    .X(_05931_));
 sky130_fd_sc_hd__nand2_1 _22010_ (.A(_05882_),
    .B(net670),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ai_1 _22011_ (.A1(_05912_),
    .A2(_05931_),
    .B1(net671),
    .Y(_01452_));
 sky130_fd_sc_hd__buf_4 _22012_ (.A(_05892_),
    .X(_05933_));
 sky130_fd_sc_hd__a211o_1 _22013_ (.A1(_05551_),
    .A2(_05884_),
    .B1(_05933_),
    .C1(_05894_),
    .X(_05934_));
 sky130_fd_sc_hd__nand2_1 _22014_ (.A(_05882_),
    .B(net1919),
    .Y(_05935_));
 sky130_fd_sc_hd__o21ai_1 _22015_ (.A1(_05912_),
    .A2(_05934_),
    .B1(net1920),
    .Y(_01453_));
 sky130_fd_sc_hd__a211o_1 _22016_ (.A1(_05555_),
    .A2(_05884_),
    .B1(_05933_),
    .C1(_05897_),
    .X(_05936_));
 sky130_fd_sc_hd__nand2_1 _22017_ (.A(_05882_),
    .B(net648),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_1 _22018_ (.A1(_05912_),
    .A2(_05936_),
    .B1(net649),
    .Y(_01454_));
 sky130_fd_sc_hd__a211o_1 _22019_ (.A1(_05558_),
    .A2(_05884_),
    .B1(_05933_),
    .C1(_05900_),
    .X(_05938_));
 sky130_fd_sc_hd__nand2_1 _22020_ (.A(_05882_),
    .B(net1929),
    .Y(_05939_));
 sky130_fd_sc_hd__o21ai_1 _22021_ (.A1(_05912_),
    .A2(_05938_),
    .B1(net1930),
    .Y(_01455_));
 sky130_fd_sc_hd__a211o_1 _22022_ (.A1(_05561_),
    .A2(_05884_),
    .B1(_05933_),
    .C1(_05903_),
    .X(_05940_));
 sky130_fd_sc_hd__nand2_1 _22023_ (.A(_05882_),
    .B(net650),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_1 _22024_ (.A1(_05912_),
    .A2(_05940_),
    .B1(net651),
    .Y(_01456_));
 sky130_fd_sc_hd__a211o_1 _22025_ (.A1(_05564_),
    .A2(_05884_),
    .B1(_05933_),
    .C1(_05906_),
    .X(_05942_));
 sky130_fd_sc_hd__nand2_1 _22026_ (.A(_05882_),
    .B(net626),
    .Y(_05943_));
 sky130_fd_sc_hd__o21ai_1 _22027_ (.A1(_05912_),
    .A2(_05942_),
    .B1(net627),
    .Y(_01457_));
 sky130_fd_sc_hd__a211o_1 _22028_ (.A1(_05567_),
    .A2(_05884_),
    .B1(_05933_),
    .C1(_05909_),
    .X(_05944_));
 sky130_fd_sc_hd__nand2_1 _22029_ (.A(_05882_),
    .B(net906),
    .Y(_05945_));
 sky130_fd_sc_hd__o21ai_1 _22030_ (.A1(_05912_),
    .A2(_05944_),
    .B1(net907),
    .Y(_01458_));
 sky130_fd_sc_hd__and3_4 _22031_ (.A(_03516_),
    .B(\line_cache_idx[7] ),
    .C(_12303_),
    .X(_05946_));
 sky130_fd_sc_hd__nand2_1 _22032_ (.A(_05946_),
    .B(_04104_),
    .Y(_05947_));
 sky130_fd_sc_hd__a21bo_1 _22033_ (.A1(_05947_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_8 _22034_ (.A(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__mux2_1 _22035_ (.A0(_05318_),
    .A1(net2298),
    .S(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__clkbuf_1 _22036_ (.A(_05950_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _22037_ (.A0(_05324_),
    .A1(net2999),
    .S(_05949_),
    .X(_05951_));
 sky130_fd_sc_hd__clkbuf_1 _22038_ (.A(_05951_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _22039_ (.A0(_05326_),
    .A1(net2505),
    .S(_05949_),
    .X(_05952_));
 sky130_fd_sc_hd__clkbuf_1 _22040_ (.A(_05952_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _22041_ (.A0(_05328_),
    .A1(net3145),
    .S(_05949_),
    .X(_05953_));
 sky130_fd_sc_hd__clkbuf_1 _22042_ (.A(_05953_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _22043_ (.A0(_05330_),
    .A1(net2603),
    .S(_05949_),
    .X(_05954_));
 sky130_fd_sc_hd__clkbuf_1 _22044_ (.A(_05954_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _22045_ (.A0(_05332_),
    .A1(net3393),
    .S(_05949_),
    .X(_05955_));
 sky130_fd_sc_hd__clkbuf_1 _22046_ (.A(_05955_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _22047_ (.A0(_05334_),
    .A1(net3422),
    .S(_05949_),
    .X(_05956_));
 sky130_fd_sc_hd__clkbuf_1 _22048_ (.A(_05956_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _22049_ (.A0(_05336_),
    .A1(net2619),
    .S(_05949_),
    .X(_05957_));
 sky130_fd_sc_hd__clkbuf_1 _22050_ (.A(_05957_),
    .X(_01466_));
 sky130_fd_sc_hd__buf_4 _22051_ (.A(_05947_),
    .X(_05958_));
 sky130_fd_sc_hd__buf_4 _22052_ (.A(_05947_),
    .X(_05959_));
 sky130_fd_sc_hd__nand2_1 _22053_ (.A(_05959_),
    .B(_05010_),
    .Y(_05960_));
 sky130_fd_sc_hd__o211a_1 _22054_ (.A1(_05095_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__mux2_1 _22055_ (.A0(_05961_),
    .A1(net2365),
    .S(_05949_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_1 _22056_ (.A(_05962_),
    .X(_01467_));
 sky130_fd_sc_hd__nand2_1 _22057_ (.A(_05959_),
    .B(_05014_),
    .Y(_05963_));
 sky130_fd_sc_hd__o211a_1 _22058_ (.A1(_05101_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__mux2_1 _22059_ (.A0(_05964_),
    .A1(net2248),
    .S(_05949_),
    .X(_05965_));
 sky130_fd_sc_hd__clkbuf_1 _22060_ (.A(_05965_),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_1 _22061_ (.A(_05959_),
    .B(_05018_),
    .Y(_05966_));
 sky130_fd_sc_hd__o211a_1 _22062_ (.A1(_05105_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__mux2_1 _22063_ (.A0(_05967_),
    .A1(net2216),
    .S(_05949_),
    .X(_05968_));
 sky130_fd_sc_hd__clkbuf_1 _22064_ (.A(_05968_),
    .X(_01469_));
 sky130_fd_sc_hd__nand2_1 _22065_ (.A(_05959_),
    .B(_05022_),
    .Y(_05969_));
 sky130_fd_sc_hd__o211a_1 _22066_ (.A1(_05109_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__mux2_1 _22067_ (.A0(_05970_),
    .A1(net2701),
    .S(_05949_),
    .X(_05971_));
 sky130_fd_sc_hd__clkbuf_1 _22068_ (.A(_05971_),
    .X(_01470_));
 sky130_fd_sc_hd__nand2_1 _22069_ (.A(_05959_),
    .B(_05026_),
    .Y(_05972_));
 sky130_fd_sc_hd__o211a_1 _22070_ (.A1(_05113_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__mux2_1 _22071_ (.A0(_05973_),
    .A1(net2539),
    .S(_05949_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _22072_ (.A(_05974_),
    .X(_01471_));
 sky130_fd_sc_hd__nand2_1 _22073_ (.A(_05959_),
    .B(_05030_),
    .Y(_05975_));
 sky130_fd_sc_hd__o211a_1 _22074_ (.A1(_05117_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__mux2_1 _22075_ (.A0(_05976_),
    .A1(net2219),
    .S(_05949_),
    .X(_05977_));
 sky130_fd_sc_hd__clkbuf_1 _22076_ (.A(_05977_),
    .X(_01472_));
 sky130_fd_sc_hd__nand2_1 _22077_ (.A(_05959_),
    .B(_05034_),
    .Y(_05978_));
 sky130_fd_sc_hd__o211a_1 _22078_ (.A1(_05121_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_1 _22079_ (.A0(_05979_),
    .A1(net2235),
    .S(_05949_),
    .X(_05980_));
 sky130_fd_sc_hd__clkbuf_1 _22080_ (.A(_05980_),
    .X(_01473_));
 sky130_fd_sc_hd__nand2_1 _22081_ (.A(_05959_),
    .B(_05038_),
    .Y(_05981_));
 sky130_fd_sc_hd__o211a_1 _22082_ (.A1(_05125_),
    .A2(_05958_),
    .B1(_05707_),
    .C1(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__mux2_1 _22083_ (.A0(_05982_),
    .A1(net3226),
    .S(_05949_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _22084_ (.A(_05983_),
    .X(_01474_));
 sky130_fd_sc_hd__buf_4 _22085_ (.A(_05183_),
    .X(_05984_));
 sky130_fd_sc_hd__o211a_1 _22086_ (.A1(_05129_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05960_),
    .X(_05985_));
 sky130_fd_sc_hd__clkbuf_8 _22087_ (.A(_05948_),
    .X(_05986_));
 sky130_fd_sc_hd__mux2_1 _22088_ (.A0(_05985_),
    .A1(net3591),
    .S(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _22089_ (.A(_05987_),
    .X(_01475_));
 sky130_fd_sc_hd__o211a_1 _22090_ (.A1(_05134_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05963_),
    .X(_05988_));
 sky130_fd_sc_hd__mux2_1 _22091_ (.A0(_05988_),
    .A1(net3461),
    .S(_05986_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_1 _22092_ (.A(_05989_),
    .X(_01476_));
 sky130_fd_sc_hd__o211a_1 _22093_ (.A1(_05137_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05966_),
    .X(_05990_));
 sky130_fd_sc_hd__mux2_1 _22094_ (.A0(_05990_),
    .A1(net3717),
    .S(_05986_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _22095_ (.A(_05991_),
    .X(_01477_));
 sky130_fd_sc_hd__o211a_1 _22096_ (.A1(_05140_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05969_),
    .X(_05992_));
 sky130_fd_sc_hd__mux2_1 _22097_ (.A0(_05992_),
    .A1(net3076),
    .S(_05986_),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_1 _22098_ (.A(_05993_),
    .X(_01478_));
 sky130_fd_sc_hd__o211a_1 _22099_ (.A1(_05143_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05972_),
    .X(_05994_));
 sky130_fd_sc_hd__mux2_1 _22100_ (.A0(_05994_),
    .A1(net3864),
    .S(_05986_),
    .X(_05995_));
 sky130_fd_sc_hd__clkbuf_1 _22101_ (.A(_05995_),
    .X(_01479_));
 sky130_fd_sc_hd__o211a_1 _22102_ (.A1(_05146_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05975_),
    .X(_05996_));
 sky130_fd_sc_hd__mux2_1 _22103_ (.A0(_05996_),
    .A1(net2230),
    .S(_05986_),
    .X(_05997_));
 sky130_fd_sc_hd__clkbuf_1 _22104_ (.A(_05997_),
    .X(_01480_));
 sky130_fd_sc_hd__o211a_1 _22105_ (.A1(_05149_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05978_),
    .X(_05998_));
 sky130_fd_sc_hd__mux2_1 _22106_ (.A0(_05998_),
    .A1(net3612),
    .S(_05986_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _22107_ (.A(_05999_),
    .X(_01481_));
 sky130_fd_sc_hd__o211a_1 _22108_ (.A1(_05152_),
    .A2(_05958_),
    .B1(_05984_),
    .C1(_05981_),
    .X(_06000_));
 sky130_fd_sc_hd__mux2_1 _22109_ (.A0(_06000_),
    .A1(net2488),
    .S(_05986_),
    .X(_06001_));
 sky130_fd_sc_hd__clkbuf_1 _22110_ (.A(_06001_),
    .X(_01482_));
 sky130_fd_sc_hd__o211a_1 _22111_ (.A1(_05059_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05960_),
    .X(_06002_));
 sky130_fd_sc_hd__mux2_1 _22112_ (.A0(_06002_),
    .A1(net3640),
    .S(_05986_),
    .X(_06003_));
 sky130_fd_sc_hd__clkbuf_1 _22113_ (.A(_06003_),
    .X(_01483_));
 sky130_fd_sc_hd__o211a_1 _22114_ (.A1(_05063_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05963_),
    .X(_06004_));
 sky130_fd_sc_hd__mux2_1 _22115_ (.A0(_06004_),
    .A1(net2047),
    .S(_05986_),
    .X(_06005_));
 sky130_fd_sc_hd__clkbuf_1 _22116_ (.A(_06005_),
    .X(_01484_));
 sky130_fd_sc_hd__o211a_1 _22117_ (.A1(_05066_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05966_),
    .X(_06006_));
 sky130_fd_sc_hd__mux2_1 _22118_ (.A0(_06006_),
    .A1(net3606),
    .S(_05986_),
    .X(_06007_));
 sky130_fd_sc_hd__clkbuf_1 _22119_ (.A(_06007_),
    .X(_01485_));
 sky130_fd_sc_hd__o211a_1 _22120_ (.A1(_05069_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05969_),
    .X(_06008_));
 sky130_fd_sc_hd__mux2_1 _22121_ (.A0(_06008_),
    .A1(net2143),
    .S(_05986_),
    .X(_06009_));
 sky130_fd_sc_hd__clkbuf_1 _22122_ (.A(_06009_),
    .X(_01486_));
 sky130_fd_sc_hd__o211a_1 _22123_ (.A1(_05072_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05972_),
    .X(_06010_));
 sky130_fd_sc_hd__mux2_1 _22124_ (.A0(_06010_),
    .A1(net3879),
    .S(_05986_),
    .X(_06011_));
 sky130_fd_sc_hd__clkbuf_1 _22125_ (.A(_06011_),
    .X(_01487_));
 sky130_fd_sc_hd__o211a_1 _22126_ (.A1(_05075_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05975_),
    .X(_06012_));
 sky130_fd_sc_hd__mux2_1 _22127_ (.A0(_06012_),
    .A1(net2256),
    .S(_05986_),
    .X(_06013_));
 sky130_fd_sc_hd__clkbuf_1 _22128_ (.A(_06013_),
    .X(_01488_));
 sky130_fd_sc_hd__o211a_1 _22129_ (.A1(_05078_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05978_),
    .X(_06014_));
 sky130_fd_sc_hd__mux2_1 _22130_ (.A0(_06014_),
    .A1(net2232),
    .S(_05986_),
    .X(_06015_));
 sky130_fd_sc_hd__clkbuf_1 _22131_ (.A(_06015_),
    .X(_01489_));
 sky130_fd_sc_hd__o211a_1 _22132_ (.A1(_05081_),
    .A2(_05959_),
    .B1(_05984_),
    .C1(_05981_),
    .X(_06016_));
 sky130_fd_sc_hd__mux2_1 _22133_ (.A0(_06016_),
    .A1(net2285),
    .S(_05986_),
    .X(_06017_));
 sky130_fd_sc_hd__clkbuf_1 _22134_ (.A(_06017_),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _22135_ (.A(_05946_),
    .B(_04183_),
    .Y(_06018_));
 sky130_fd_sc_hd__inv_2 _22136_ (.A(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__clkbuf_16 _22137_ (.A(_12190_),
    .X(_06020_));
 sky130_fd_sc_hd__o21ai_4 _22138_ (.A1(_05471_),
    .A2(_06019_),
    .B1(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__mux2_1 _22139_ (.A0(_05318_),
    .A1(net3559),
    .S(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__clkbuf_1 _22140_ (.A(_06022_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _22141_ (.A0(_05324_),
    .A1(net3628),
    .S(_06021_),
    .X(_06023_));
 sky130_fd_sc_hd__clkbuf_1 _22142_ (.A(_06023_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _22143_ (.A0(_05326_),
    .A1(net3269),
    .S(_06021_),
    .X(_06024_));
 sky130_fd_sc_hd__clkbuf_1 _22144_ (.A(_06024_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _22145_ (.A0(_05328_),
    .A1(net3255),
    .S(_06021_),
    .X(_06025_));
 sky130_fd_sc_hd__clkbuf_1 _22146_ (.A(_06025_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _22147_ (.A0(_05330_),
    .A1(net2695),
    .S(_06021_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _22148_ (.A(_06026_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _22149_ (.A0(_05332_),
    .A1(net3302),
    .S(_06021_),
    .X(_06027_));
 sky130_fd_sc_hd__clkbuf_1 _22150_ (.A(_06027_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _22151_ (.A0(_05334_),
    .A1(net3682),
    .S(_06021_),
    .X(_06028_));
 sky130_fd_sc_hd__clkbuf_1 _22152_ (.A(_06028_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _22153_ (.A0(_05336_),
    .A1(net3324),
    .S(_06021_),
    .X(_06029_));
 sky130_fd_sc_hd__clkbuf_1 _22154_ (.A(_06029_),
    .X(_01498_));
 sky130_fd_sc_hd__buf_4 _22155_ (.A(_06021_),
    .X(_06030_));
 sky130_fd_sc_hd__buf_4 _22156_ (.A(_06019_),
    .X(_06031_));
 sky130_fd_sc_hd__buf_4 _22157_ (.A(_06019_),
    .X(_06032_));
 sky130_fd_sc_hd__nor2_1 _22158_ (.A(_05583_),
    .B(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__a211o_1 _22159_ (.A1(_05484_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__buf_4 _22160_ (.A(_06021_),
    .X(_06035_));
 sky130_fd_sc_hd__nand2_1 _22161_ (.A(_06035_),
    .B(net1036),
    .Y(_06036_));
 sky130_fd_sc_hd__o21ai_1 _22162_ (.A1(_06030_),
    .A2(_06034_),
    .B1(net1037),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_05589_),
    .B(_06032_),
    .Y(_06037_));
 sky130_fd_sc_hd__a211o_1 _22164_ (.A1(_05491_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__nand2_1 _22165_ (.A(_06035_),
    .B(net1398),
    .Y(_06039_));
 sky130_fd_sc_hd__o21ai_1 _22166_ (.A1(_06030_),
    .A2(_06038_),
    .B1(net1399),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _22167_ (.A(_05593_),
    .B(_06032_),
    .Y(_06040_));
 sky130_fd_sc_hd__a211o_1 _22168_ (.A1(_05495_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2_1 _22169_ (.A(_06035_),
    .B(net1506),
    .Y(_06042_));
 sky130_fd_sc_hd__o21ai_1 _22170_ (.A1(_06030_),
    .A2(_06041_),
    .B1(net1507),
    .Y(_01501_));
 sky130_fd_sc_hd__nor2_1 _22171_ (.A(_05597_),
    .B(_06032_),
    .Y(_06043_));
 sky130_fd_sc_hd__a211o_1 _22172_ (.A1(_05500_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__nand2_1 _22173_ (.A(_06035_),
    .B(net1804),
    .Y(_06045_));
 sky130_fd_sc_hd__o21ai_1 _22174_ (.A1(_06030_),
    .A2(_06044_),
    .B1(net1805),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _22175_ (.A(_05601_),
    .B(_06032_),
    .Y(_06046_));
 sky130_fd_sc_hd__a211o_1 _22176_ (.A1(_05504_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__nand2_1 _22177_ (.A(_06035_),
    .B(net1022),
    .Y(_06048_));
 sky130_fd_sc_hd__o21ai_1 _22178_ (.A1(_06030_),
    .A2(_06047_),
    .B1(net1023),
    .Y(_01503_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_05605_),
    .B(_06032_),
    .Y(_06049_));
 sky130_fd_sc_hd__a211o_1 _22180_ (.A1(_05508_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__nand2_1 _22181_ (.A(_06035_),
    .B(net1518),
    .Y(_06051_));
 sky130_fd_sc_hd__o21ai_1 _22182_ (.A1(_06030_),
    .A2(_06050_),
    .B1(net1519),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_1 _22183_ (.A(_05609_),
    .B(_06032_),
    .Y(_06052_));
 sky130_fd_sc_hd__a211o_1 _22184_ (.A1(_05512_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__nand2_1 _22185_ (.A(_06035_),
    .B(net1340),
    .Y(_06054_));
 sky130_fd_sc_hd__o21ai_1 _22186_ (.A1(_06030_),
    .A2(_06053_),
    .B1(net1341),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _22187_ (.A(_05613_),
    .B(_06032_),
    .Y(_06055_));
 sky130_fd_sc_hd__a211o_1 _22188_ (.A1(_05516_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__nand2_1 _22189_ (.A(_06035_),
    .B(net1214),
    .Y(_06057_));
 sky130_fd_sc_hd__o21ai_1 _22190_ (.A1(_06030_),
    .A2(_06056_),
    .B1(net1215),
    .Y(_01506_));
 sky130_fd_sc_hd__buf_4 _22191_ (.A(_06021_),
    .X(_06058_));
 sky130_fd_sc_hd__a211o_1 _22192_ (.A1(_05521_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06033_),
    .X(_06059_));
 sky130_fd_sc_hd__nand2_1 _22193_ (.A(_06035_),
    .B(net1354),
    .Y(_06060_));
 sky130_fd_sc_hd__o21ai_1 _22194_ (.A1(_06058_),
    .A2(_06059_),
    .B1(net1355),
    .Y(_01507_));
 sky130_fd_sc_hd__a211o_1 _22195_ (.A1(_05524_),
    .A2(_06031_),
    .B1(_05933_),
    .C1(_06037_),
    .X(_06061_));
 sky130_fd_sc_hd__nand2_1 _22196_ (.A(_06035_),
    .B(net1676),
    .Y(_06062_));
 sky130_fd_sc_hd__o21ai_1 _22197_ (.A1(_06058_),
    .A2(_06061_),
    .B1(net1677),
    .Y(_01508_));
 sky130_fd_sc_hd__buf_4 _22198_ (.A(_05892_),
    .X(_06063_));
 sky130_fd_sc_hd__a211o_1 _22199_ (.A1(_05527_),
    .A2(_06031_),
    .B1(_06063_),
    .C1(_06040_),
    .X(_06064_));
 sky130_fd_sc_hd__nand2_1 _22200_ (.A(_06035_),
    .B(net538),
    .Y(_06065_));
 sky130_fd_sc_hd__o21ai_1 _22201_ (.A1(_06058_),
    .A2(_06064_),
    .B1(net539),
    .Y(_01509_));
 sky130_fd_sc_hd__a211o_1 _22202_ (.A1(_05530_),
    .A2(_06031_),
    .B1(_06063_),
    .C1(_06043_),
    .X(_06066_));
 sky130_fd_sc_hd__nand2_1 _22203_ (.A(_06035_),
    .B(net1090),
    .Y(_06067_));
 sky130_fd_sc_hd__o21ai_1 _22204_ (.A1(_06058_),
    .A2(_06066_),
    .B1(net1091),
    .Y(_01510_));
 sky130_fd_sc_hd__a211o_1 _22205_ (.A1(_05533_),
    .A2(_06031_),
    .B1(_06063_),
    .C1(_06046_),
    .X(_06068_));
 sky130_fd_sc_hd__nand2_1 _22206_ (.A(_06035_),
    .B(net804),
    .Y(_06069_));
 sky130_fd_sc_hd__o21ai_1 _22207_ (.A1(_06058_),
    .A2(_06068_),
    .B1(net805),
    .Y(_01511_));
 sky130_fd_sc_hd__a211o_1 _22208_ (.A1(_05536_),
    .A2(_06031_),
    .B1(_06063_),
    .C1(_06049_),
    .X(_06070_));
 sky130_fd_sc_hd__nand2_1 _22209_ (.A(_06035_),
    .B(net1444),
    .Y(_06071_));
 sky130_fd_sc_hd__o21ai_1 _22210_ (.A1(_06058_),
    .A2(_06070_),
    .B1(net1445),
    .Y(_01512_));
 sky130_fd_sc_hd__a211o_1 _22211_ (.A1(_05539_),
    .A2(_06031_),
    .B1(_06063_),
    .C1(_06052_),
    .X(_06072_));
 sky130_fd_sc_hd__nand2_1 _22212_ (.A(_06035_),
    .B(net1460),
    .Y(_06073_));
 sky130_fd_sc_hd__o21ai_1 _22213_ (.A1(_06058_),
    .A2(_06072_),
    .B1(net1461),
    .Y(_01513_));
 sky130_fd_sc_hd__a211o_1 _22214_ (.A1(_05542_),
    .A2(_06031_),
    .B1(_06063_),
    .C1(_06055_),
    .X(_06074_));
 sky130_fd_sc_hd__nand2_1 _22215_ (.A(_06035_),
    .B(net1386),
    .Y(_06075_));
 sky130_fd_sc_hd__o21ai_1 _22216_ (.A1(_06058_),
    .A2(_06074_),
    .B1(net1387),
    .Y(_01514_));
 sky130_fd_sc_hd__a211o_1 _22217_ (.A1(_05545_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06033_),
    .X(_06076_));
 sky130_fd_sc_hd__nand2_1 _22218_ (.A(_06030_),
    .B(net1366),
    .Y(_06077_));
 sky130_fd_sc_hd__o21ai_1 _22219_ (.A1(_06058_),
    .A2(_06076_),
    .B1(net1367),
    .Y(_01515_));
 sky130_fd_sc_hd__a211o_1 _22220_ (.A1(_05548_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06037_),
    .X(_06078_));
 sky130_fd_sc_hd__nand2_1 _22221_ (.A(_06030_),
    .B(net684),
    .Y(_06079_));
 sky130_fd_sc_hd__o21ai_1 _22222_ (.A1(_06058_),
    .A2(_06078_),
    .B1(net685),
    .Y(_01516_));
 sky130_fd_sc_hd__a211o_1 _22223_ (.A1(_05551_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06040_),
    .X(_06080_));
 sky130_fd_sc_hd__nand2_1 _22224_ (.A(_06030_),
    .B(net1724),
    .Y(_06081_));
 sky130_fd_sc_hd__o21ai_1 _22225_ (.A1(_06058_),
    .A2(_06080_),
    .B1(net1725),
    .Y(_01517_));
 sky130_fd_sc_hd__a211o_1 _22226_ (.A1(_05555_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06043_),
    .X(_06082_));
 sky130_fd_sc_hd__nand2_1 _22227_ (.A(_06030_),
    .B(net1788),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_1 _22228_ (.A1(_06058_),
    .A2(_06082_),
    .B1(net1789),
    .Y(_01518_));
 sky130_fd_sc_hd__a211o_1 _22229_ (.A1(_05558_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06046_),
    .X(_06084_));
 sky130_fd_sc_hd__nand2_1 _22230_ (.A(_06030_),
    .B(net1838),
    .Y(_06085_));
 sky130_fd_sc_hd__o21ai_1 _22231_ (.A1(_06058_),
    .A2(_06084_),
    .B1(net1839),
    .Y(_01519_));
 sky130_fd_sc_hd__a211o_1 _22232_ (.A1(_05561_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06049_),
    .X(_06086_));
 sky130_fd_sc_hd__nand2_1 _22233_ (.A(_06030_),
    .B(net1856),
    .Y(_06087_));
 sky130_fd_sc_hd__o21ai_1 _22234_ (.A1(_06058_),
    .A2(_06086_),
    .B1(net1857),
    .Y(_01520_));
 sky130_fd_sc_hd__a211o_1 _22235_ (.A1(_05564_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06052_),
    .X(_06088_));
 sky130_fd_sc_hd__nand2_1 _22236_ (.A(_06030_),
    .B(net644),
    .Y(_06089_));
 sky130_fd_sc_hd__o21ai_1 _22237_ (.A1(_06058_),
    .A2(_06088_),
    .B1(net645),
    .Y(_01521_));
 sky130_fd_sc_hd__a211o_1 _22238_ (.A1(_05567_),
    .A2(_06032_),
    .B1(_06063_),
    .C1(_06055_),
    .X(_06090_));
 sky130_fd_sc_hd__nand2_1 _22239_ (.A(_06030_),
    .B(net1642),
    .Y(_06091_));
 sky130_fd_sc_hd__o21ai_1 _22240_ (.A1(_06058_),
    .A2(_06090_),
    .B1(net1643),
    .Y(_01522_));
 sky130_fd_sc_hd__nand2_1 _22241_ (.A(_05946_),
    .B(_04257_),
    .Y(_06092_));
 sky130_fd_sc_hd__inv_2 _22242_ (.A(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__o21ai_4 _22243_ (.A1(_05471_),
    .A2(_06093_),
    .B1(_06020_),
    .Y(_06094_));
 sky130_fd_sc_hd__mux2_1 _22244_ (.A0(_05318_),
    .A1(net3719),
    .S(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__clkbuf_1 _22245_ (.A(_06095_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _22246_ (.A0(_05324_),
    .A1(net2835),
    .S(_06094_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _22247_ (.A(_06096_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _22248_ (.A0(_05326_),
    .A1(net3057),
    .S(_06094_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _22249_ (.A(_06097_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _22250_ (.A0(_05328_),
    .A1(net2770),
    .S(_06094_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _22251_ (.A(_06098_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _22252_ (.A0(_05330_),
    .A1(net2785),
    .S(_06094_),
    .X(_06099_));
 sky130_fd_sc_hd__clkbuf_1 _22253_ (.A(_06099_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _22254_ (.A0(_05332_),
    .A1(net2906),
    .S(_06094_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_1 _22255_ (.A(_06100_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _22256_ (.A0(_05334_),
    .A1(net3314),
    .S(_06094_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _22257_ (.A(_06101_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _22258_ (.A0(_05336_),
    .A1(net2852),
    .S(_06094_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_1 _22259_ (.A(_06102_),
    .X(_01530_));
 sky130_fd_sc_hd__buf_4 _22260_ (.A(_06094_),
    .X(_06103_));
 sky130_fd_sc_hd__buf_4 _22261_ (.A(_06093_),
    .X(_06104_));
 sky130_fd_sc_hd__buf_4 _22262_ (.A(_06093_),
    .X(_06105_));
 sky130_fd_sc_hd__nor2_1 _22263_ (.A(_05583_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__a211o_1 _22264_ (.A1(_05484_),
    .A2(_06104_),
    .B1(_06063_),
    .C1(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__buf_4 _22265_ (.A(_06094_),
    .X(_06108_));
 sky130_fd_sc_hd__nand2_1 _22266_ (.A(_06108_),
    .B(net1954),
    .Y(_06109_));
 sky130_fd_sc_hd__o21ai_1 _22267_ (.A1(_06103_),
    .A2(_06107_),
    .B1(_06109_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _22268_ (.A(_05589_),
    .B(_06105_),
    .Y(_06110_));
 sky130_fd_sc_hd__a211o_1 _22269_ (.A1(_05491_),
    .A2(_06104_),
    .B1(_06063_),
    .C1(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__nand2_1 _22270_ (.A(_06108_),
    .B(net1126),
    .Y(_06112_));
 sky130_fd_sc_hd__o21ai_1 _22271_ (.A1(_06103_),
    .A2(_06111_),
    .B1(net1127),
    .Y(_01532_));
 sky130_fd_sc_hd__buf_4 _22272_ (.A(_05892_),
    .X(_06113_));
 sky130_fd_sc_hd__nor2_1 _22273_ (.A(_05593_),
    .B(_06105_),
    .Y(_06114_));
 sky130_fd_sc_hd__a211o_1 _22274_ (.A1(_05495_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__nand2_1 _22275_ (.A(_06108_),
    .B(net980),
    .Y(_06116_));
 sky130_fd_sc_hd__o21ai_1 _22276_ (.A1(_06103_),
    .A2(_06115_),
    .B1(net981),
    .Y(_01533_));
 sky130_fd_sc_hd__nor2_1 _22277_ (.A(_05597_),
    .B(_06105_),
    .Y(_06117_));
 sky130_fd_sc_hd__a211o_1 _22278_ (.A1(_05500_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__nand2_1 _22279_ (.A(_06108_),
    .B(net1094),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_1 _22280_ (.A1(_06103_),
    .A2(_06118_),
    .B1(net1095),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _22281_ (.A(_05601_),
    .B(_06105_),
    .Y(_06120_));
 sky130_fd_sc_hd__a211o_1 _22282_ (.A1(_05504_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__nand2_1 _22283_ (.A(_06108_),
    .B(net880),
    .Y(_06122_));
 sky130_fd_sc_hd__o21ai_1 _22284_ (.A1(_06103_),
    .A2(_06121_),
    .B1(net881),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _22285_ (.A(_05605_),
    .B(_06105_),
    .Y(_06123_));
 sky130_fd_sc_hd__a211o_1 _22286_ (.A1(_05508_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__nand2_1 _22287_ (.A(_06108_),
    .B(net1486),
    .Y(_06125_));
 sky130_fd_sc_hd__o21ai_1 _22288_ (.A1(_06103_),
    .A2(_06124_),
    .B1(net1487),
    .Y(_01536_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(_05609_),
    .B(_06105_),
    .Y(_06126_));
 sky130_fd_sc_hd__a211o_1 _22290_ (.A1(_05512_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06126_),
    .X(_06127_));
 sky130_fd_sc_hd__nand2_1 _22291_ (.A(_06108_),
    .B(net1060),
    .Y(_06128_));
 sky130_fd_sc_hd__o21ai_1 _22292_ (.A1(_06103_),
    .A2(_06127_),
    .B1(net1061),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _22293_ (.A(_05613_),
    .B(_06105_),
    .Y(_06129_));
 sky130_fd_sc_hd__a211o_1 _22294_ (.A1(_05516_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__nand2_1 _22295_ (.A(_06108_),
    .B(net564),
    .Y(_06131_));
 sky130_fd_sc_hd__o21ai_1 _22296_ (.A1(_06103_),
    .A2(_06130_),
    .B1(net565),
    .Y(_01538_));
 sky130_fd_sc_hd__buf_4 _22297_ (.A(_06094_),
    .X(_06132_));
 sky130_fd_sc_hd__a211o_1 _22298_ (.A1(_05521_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06106_),
    .X(_06133_));
 sky130_fd_sc_hd__nand2_1 _22299_ (.A(_06108_),
    .B(net1678),
    .Y(_06134_));
 sky130_fd_sc_hd__o21ai_1 _22300_ (.A1(_06132_),
    .A2(_06133_),
    .B1(net1679),
    .Y(_01539_));
 sky130_fd_sc_hd__a211o_1 _22301_ (.A1(_05524_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06110_),
    .X(_06135_));
 sky130_fd_sc_hd__nand2_1 _22302_ (.A(_06108_),
    .B(net1068),
    .Y(_06136_));
 sky130_fd_sc_hd__o21ai_1 _22303_ (.A1(_06132_),
    .A2(_06135_),
    .B1(net1069),
    .Y(_01540_));
 sky130_fd_sc_hd__a211o_1 _22304_ (.A1(_05527_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06114_),
    .X(_06137_));
 sky130_fd_sc_hd__nand2_1 _22305_ (.A(_06108_),
    .B(net1943),
    .Y(_06138_));
 sky130_fd_sc_hd__o21ai_1 _22306_ (.A1(_06132_),
    .A2(_06137_),
    .B1(_06138_),
    .Y(_01541_));
 sky130_fd_sc_hd__a211o_1 _22307_ (.A1(_05530_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06117_),
    .X(_06139_));
 sky130_fd_sc_hd__nand2_1 _22308_ (.A(_06108_),
    .B(net920),
    .Y(_06140_));
 sky130_fd_sc_hd__o21ai_1 _22309_ (.A1(_06132_),
    .A2(_06139_),
    .B1(net921),
    .Y(_01542_));
 sky130_fd_sc_hd__a211o_1 _22310_ (.A1(_05533_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06120_),
    .X(_06141_));
 sky130_fd_sc_hd__nand2_1 _22311_ (.A(_06108_),
    .B(net1966),
    .Y(_06142_));
 sky130_fd_sc_hd__o21ai_1 _22312_ (.A1(_06132_),
    .A2(_06141_),
    .B1(_06142_),
    .Y(_01543_));
 sky130_fd_sc_hd__a211o_1 _22313_ (.A1(_05536_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06123_),
    .X(_06143_));
 sky130_fd_sc_hd__nand2_1 _22314_ (.A(_06108_),
    .B(net1630),
    .Y(_06144_));
 sky130_fd_sc_hd__o21ai_1 _22315_ (.A1(_06132_),
    .A2(_06143_),
    .B1(net1631),
    .Y(_01544_));
 sky130_fd_sc_hd__a211o_1 _22316_ (.A1(_05539_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06126_),
    .X(_06145_));
 sky130_fd_sc_hd__nand2_1 _22317_ (.A(_06108_),
    .B(net1406),
    .Y(_06146_));
 sky130_fd_sc_hd__o21ai_1 _22318_ (.A1(_06132_),
    .A2(_06145_),
    .B1(net1407),
    .Y(_01545_));
 sky130_fd_sc_hd__a211o_1 _22319_ (.A1(_05542_),
    .A2(_06104_),
    .B1(_06113_),
    .C1(_06129_),
    .X(_06147_));
 sky130_fd_sc_hd__nand2_1 _22320_ (.A(_06108_),
    .B(net1322),
    .Y(_06148_));
 sky130_fd_sc_hd__o21ai_1 _22321_ (.A1(_06132_),
    .A2(_06147_),
    .B1(net1323),
    .Y(_01546_));
 sky130_fd_sc_hd__a211o_1 _22322_ (.A1(_05545_),
    .A2(_06105_),
    .B1(_06113_),
    .C1(_06106_),
    .X(_06149_));
 sky130_fd_sc_hd__nand2_1 _22323_ (.A(_06103_),
    .B(net1462),
    .Y(_06150_));
 sky130_fd_sc_hd__o21ai_1 _22324_ (.A1(_06132_),
    .A2(_06149_),
    .B1(net1463),
    .Y(_01547_));
 sky130_fd_sc_hd__a211o_1 _22325_ (.A1(_05548_),
    .A2(_06105_),
    .B1(_06113_),
    .C1(_06110_),
    .X(_06151_));
 sky130_fd_sc_hd__nand2_1 _22326_ (.A(_06103_),
    .B(net1174),
    .Y(_06152_));
 sky130_fd_sc_hd__o21ai_1 _22327_ (.A1(_06132_),
    .A2(_06151_),
    .B1(net1175),
    .Y(_01548_));
 sky130_fd_sc_hd__buf_4 _22328_ (.A(_05892_),
    .X(_06153_));
 sky130_fd_sc_hd__a211o_1 _22329_ (.A1(_05551_),
    .A2(_06105_),
    .B1(_06153_),
    .C1(_06114_),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_1 _22330_ (.A(_06103_),
    .B(net1952),
    .Y(_06155_));
 sky130_fd_sc_hd__o21ai_1 _22331_ (.A1(_06132_),
    .A2(_06154_),
    .B1(_06155_),
    .Y(_01549_));
 sky130_fd_sc_hd__a211o_1 _22332_ (.A1(_05555_),
    .A2(_06105_),
    .B1(_06153_),
    .C1(_06117_),
    .X(_06156_));
 sky130_fd_sc_hd__nand2_1 _22333_ (.A(_06103_),
    .B(net574),
    .Y(_06157_));
 sky130_fd_sc_hd__o21ai_1 _22334_ (.A1(_06132_),
    .A2(_06156_),
    .B1(net575),
    .Y(_01550_));
 sky130_fd_sc_hd__a211o_1 _22335_ (.A1(_05558_),
    .A2(_06105_),
    .B1(_06153_),
    .C1(_06120_),
    .X(_06158_));
 sky130_fd_sc_hd__nand2_1 _22336_ (.A(_06103_),
    .B(net1964),
    .Y(_06159_));
 sky130_fd_sc_hd__o21ai_1 _22337_ (.A1(_06132_),
    .A2(_06158_),
    .B1(net1965),
    .Y(_01551_));
 sky130_fd_sc_hd__a211o_1 _22338_ (.A1(_05561_),
    .A2(_06105_),
    .B1(_06153_),
    .C1(_06123_),
    .X(_06160_));
 sky130_fd_sc_hd__nand2_1 _22339_ (.A(_06103_),
    .B(net1652),
    .Y(_06161_));
 sky130_fd_sc_hd__o21ai_1 _22340_ (.A1(_06132_),
    .A2(_06160_),
    .B1(net1653),
    .Y(_01552_));
 sky130_fd_sc_hd__a211o_1 _22341_ (.A1(_05564_),
    .A2(_06105_),
    .B1(_06153_),
    .C1(_06126_),
    .X(_06162_));
 sky130_fd_sc_hd__nand2_1 _22342_ (.A(_06103_),
    .B(net1070),
    .Y(_06163_));
 sky130_fd_sc_hd__o21ai_1 _22343_ (.A1(_06132_),
    .A2(_06162_),
    .B1(net1071),
    .Y(_01553_));
 sky130_fd_sc_hd__a211o_1 _22344_ (.A1(_05567_),
    .A2(_06105_),
    .B1(_06153_),
    .C1(_06129_),
    .X(_06164_));
 sky130_fd_sc_hd__nand2_1 _22345_ (.A(_06103_),
    .B(net824),
    .Y(_06165_));
 sky130_fd_sc_hd__o21ai_1 _22346_ (.A1(_06132_),
    .A2(_06164_),
    .B1(net825),
    .Y(_01554_));
 sky130_fd_sc_hd__nand2_1 _22347_ (.A(_05946_),
    .B(_04333_),
    .Y(_06166_));
 sky130_fd_sc_hd__inv_2 _22348_ (.A(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__o21ai_4 _22349_ (.A1(_05471_),
    .A2(_06167_),
    .B1(_06020_),
    .Y(_06168_));
 sky130_fd_sc_hd__mux2_1 _22350_ (.A0(_05318_),
    .A1(net3443),
    .S(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_1 _22351_ (.A(_06169_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _22352_ (.A0(_05324_),
    .A1(net3260),
    .S(_06168_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _22353_ (.A(_06170_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _22354_ (.A0(_05326_),
    .A1(net3428),
    .S(_06168_),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _22355_ (.A(_06171_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _22356_ (.A0(_05328_),
    .A1(net3809),
    .S(_06168_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _22357_ (.A(_06172_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _22358_ (.A0(_05330_),
    .A1(net2778),
    .S(_06168_),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _22359_ (.A(_06173_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _22360_ (.A0(_05332_),
    .A1(net2565),
    .S(_06168_),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _22361_ (.A(_06174_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _22362_ (.A0(_05334_),
    .A1(net3583),
    .S(_06168_),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_1 _22363_ (.A(_06175_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _22364_ (.A0(_05336_),
    .A1(net3710),
    .S(_06168_),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _22365_ (.A(_06176_),
    .X(_01562_));
 sky130_fd_sc_hd__buf_4 _22366_ (.A(_06168_),
    .X(_06177_));
 sky130_fd_sc_hd__buf_4 _22367_ (.A(_06167_),
    .X(_06178_));
 sky130_fd_sc_hd__buf_4 _22368_ (.A(_06167_),
    .X(_06179_));
 sky130_fd_sc_hd__nor2_1 _22369_ (.A(_05583_),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__a211o_1 _22370_ (.A1(_05484_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__buf_4 _22371_ (.A(_06168_),
    .X(_06182_));
 sky130_fd_sc_hd__nand2_1 _22372_ (.A(_06182_),
    .B(net1458),
    .Y(_06183_));
 sky130_fd_sc_hd__o21ai_1 _22373_ (.A1(_06177_),
    .A2(_06181_),
    .B1(net1459),
    .Y(_01563_));
 sky130_fd_sc_hd__nor2_1 _22374_ (.A(_05589_),
    .B(_06179_),
    .Y(_06184_));
 sky130_fd_sc_hd__a211o_1 _22375_ (.A1(_05491_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__nand2_1 _22376_ (.A(_06182_),
    .B(net1196),
    .Y(_06186_));
 sky130_fd_sc_hd__o21ai_1 _22377_ (.A1(_06177_),
    .A2(_06185_),
    .B1(net1197),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _22378_ (.A(_05593_),
    .B(_06179_),
    .Y(_06187_));
 sky130_fd_sc_hd__a211o_1 _22379_ (.A1(_05495_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__nand2_1 _22380_ (.A(_06182_),
    .B(net1028),
    .Y(_06189_));
 sky130_fd_sc_hd__o21ai_1 _22381_ (.A1(_06177_),
    .A2(_06188_),
    .B1(net1029),
    .Y(_01565_));
 sky130_fd_sc_hd__nor2_1 _22382_ (.A(_05597_),
    .B(_06179_),
    .Y(_06190_));
 sky130_fd_sc_hd__a211o_1 _22383_ (.A1(_05500_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__nand2_1 _22384_ (.A(_06182_),
    .B(net1058),
    .Y(_06192_));
 sky130_fd_sc_hd__o21ai_1 _22385_ (.A1(_06177_),
    .A2(_06191_),
    .B1(net1059),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _22386_ (.A(_05601_),
    .B(_06179_),
    .Y(_06193_));
 sky130_fd_sc_hd__a211o_1 _22387_ (.A1(_05504_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__nand2_1 _22388_ (.A(_06182_),
    .B(net1456),
    .Y(_06195_));
 sky130_fd_sc_hd__o21ai_1 _22389_ (.A1(_06177_),
    .A2(_06194_),
    .B1(net1457),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_1 _22390_ (.A(_05605_),
    .B(_06179_),
    .Y(_06196_));
 sky130_fd_sc_hd__a211o_1 _22391_ (.A1(_05508_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__nand2_1 _22392_ (.A(_06182_),
    .B(net1312),
    .Y(_06198_));
 sky130_fd_sc_hd__o21ai_1 _22393_ (.A1(_06177_),
    .A2(_06197_),
    .B1(net1313),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_1 _22394_ (.A(_05609_),
    .B(_06179_),
    .Y(_06199_));
 sky130_fd_sc_hd__a211o_1 _22395_ (.A1(_05512_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__nand2_1 _22396_ (.A(_06182_),
    .B(net1648),
    .Y(_06201_));
 sky130_fd_sc_hd__o21ai_1 _22397_ (.A1(_06177_),
    .A2(_06200_),
    .B1(net1649),
    .Y(_01569_));
 sky130_fd_sc_hd__nor2_1 _22398_ (.A(_05613_),
    .B(_06179_),
    .Y(_06202_));
 sky130_fd_sc_hd__a211o_1 _22399_ (.A1(_05516_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__nand2_1 _22400_ (.A(_06182_),
    .B(net986),
    .Y(_06204_));
 sky130_fd_sc_hd__o21ai_1 _22401_ (.A1(_06177_),
    .A2(_06203_),
    .B1(net987),
    .Y(_01570_));
 sky130_fd_sc_hd__buf_4 _22402_ (.A(_06168_),
    .X(_06205_));
 sky130_fd_sc_hd__a211o_1 _22403_ (.A1(_05521_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06180_),
    .X(_06206_));
 sky130_fd_sc_hd__nand2_1 _22404_ (.A(_06182_),
    .B(net994),
    .Y(_06207_));
 sky130_fd_sc_hd__o21ai_1 _22405_ (.A1(_06205_),
    .A2(_06206_),
    .B1(net995),
    .Y(_01571_));
 sky130_fd_sc_hd__a211o_1 _22406_ (.A1(_05524_),
    .A2(_06178_),
    .B1(_06153_),
    .C1(_06184_),
    .X(_06208_));
 sky130_fd_sc_hd__nand2_1 _22407_ (.A(_06182_),
    .B(net836),
    .Y(_06209_));
 sky130_fd_sc_hd__o21ai_1 _22408_ (.A1(_06205_),
    .A2(_06208_),
    .B1(net837),
    .Y(_01572_));
 sky130_fd_sc_hd__buf_4 _22409_ (.A(_05892_),
    .X(_06210_));
 sky130_fd_sc_hd__a211o_1 _22410_ (.A1(_05527_),
    .A2(_06178_),
    .B1(_06210_),
    .C1(_06187_),
    .X(_06211_));
 sky130_fd_sc_hd__nand2_1 _22411_ (.A(_06182_),
    .B(net576),
    .Y(_06212_));
 sky130_fd_sc_hd__o21ai_1 _22412_ (.A1(_06205_),
    .A2(_06211_),
    .B1(net577),
    .Y(_01573_));
 sky130_fd_sc_hd__a211o_1 _22413_ (.A1(_05530_),
    .A2(_06178_),
    .B1(_06210_),
    .C1(_06190_),
    .X(_06213_));
 sky130_fd_sc_hd__nand2_1 _22414_ (.A(_06182_),
    .B(net1598),
    .Y(_06214_));
 sky130_fd_sc_hd__o21ai_1 _22415_ (.A1(_06205_),
    .A2(_06213_),
    .B1(net1599),
    .Y(_01574_));
 sky130_fd_sc_hd__a211o_1 _22416_ (.A1(_05533_),
    .A2(_06178_),
    .B1(_06210_),
    .C1(_06193_),
    .X(_06215_));
 sky130_fd_sc_hd__nand2_1 _22417_ (.A(_06182_),
    .B(net1180),
    .Y(_06216_));
 sky130_fd_sc_hd__o21ai_1 _22418_ (.A1(_06205_),
    .A2(_06215_),
    .B1(net1181),
    .Y(_01575_));
 sky130_fd_sc_hd__a211o_1 _22419_ (.A1(_05536_),
    .A2(_06178_),
    .B1(_06210_),
    .C1(_06196_),
    .X(_06217_));
 sky130_fd_sc_hd__nand2_1 _22420_ (.A(_06182_),
    .B(net846),
    .Y(_06218_));
 sky130_fd_sc_hd__o21ai_1 _22421_ (.A1(_06205_),
    .A2(_06217_),
    .B1(net847),
    .Y(_01576_));
 sky130_fd_sc_hd__a211o_1 _22422_ (.A1(_05539_),
    .A2(_06178_),
    .B1(_06210_),
    .C1(_06199_),
    .X(_06219_));
 sky130_fd_sc_hd__nand2_1 _22423_ (.A(_06182_),
    .B(net1194),
    .Y(_06220_));
 sky130_fd_sc_hd__o21ai_1 _22424_ (.A1(_06205_),
    .A2(_06219_),
    .B1(net1195),
    .Y(_01577_));
 sky130_fd_sc_hd__a211o_1 _22425_ (.A1(_05542_),
    .A2(_06178_),
    .B1(_06210_),
    .C1(_06202_),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _22426_ (.A(_06182_),
    .B(net800),
    .Y(_06222_));
 sky130_fd_sc_hd__o21ai_1 _22427_ (.A1(_06205_),
    .A2(_06221_),
    .B1(net801),
    .Y(_01578_));
 sky130_fd_sc_hd__a211o_1 _22428_ (.A1(_05545_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06180_),
    .X(_06223_));
 sky130_fd_sc_hd__nand2_1 _22429_ (.A(_06177_),
    .B(net898),
    .Y(_06224_));
 sky130_fd_sc_hd__o21ai_1 _22430_ (.A1(_06205_),
    .A2(_06223_),
    .B1(net899),
    .Y(_01579_));
 sky130_fd_sc_hd__a211o_1 _22431_ (.A1(_05548_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06184_),
    .X(_06225_));
 sky130_fd_sc_hd__nand2_1 _22432_ (.A(_06177_),
    .B(net722),
    .Y(_06226_));
 sky130_fd_sc_hd__o21ai_1 _22433_ (.A1(_06205_),
    .A2(_06225_),
    .B1(net723),
    .Y(_01580_));
 sky130_fd_sc_hd__a211o_1 _22434_ (.A1(_05551_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06187_),
    .X(_06227_));
 sky130_fd_sc_hd__nand2_1 _22435_ (.A(_06177_),
    .B(net938),
    .Y(_06228_));
 sky130_fd_sc_hd__o21ai_1 _22436_ (.A1(_06205_),
    .A2(_06227_),
    .B1(net939),
    .Y(_01581_));
 sky130_fd_sc_hd__a211o_1 _22437_ (.A1(_05555_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06190_),
    .X(_06229_));
 sky130_fd_sc_hd__nand2_1 _22438_ (.A(_06177_),
    .B(net1358),
    .Y(_06230_));
 sky130_fd_sc_hd__o21ai_1 _22439_ (.A1(_06205_),
    .A2(_06229_),
    .B1(net1359),
    .Y(_01582_));
 sky130_fd_sc_hd__a211o_1 _22440_ (.A1(_05558_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06193_),
    .X(_06231_));
 sky130_fd_sc_hd__nand2_1 _22441_ (.A(_06177_),
    .B(net1096),
    .Y(_06232_));
 sky130_fd_sc_hd__o21ai_1 _22442_ (.A1(_06205_),
    .A2(_06231_),
    .B1(net1097),
    .Y(_01583_));
 sky130_fd_sc_hd__a211o_1 _22443_ (.A1(_05561_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06196_),
    .X(_06233_));
 sky130_fd_sc_hd__nand2_1 _22444_ (.A(_06177_),
    .B(net1632),
    .Y(_06234_));
 sky130_fd_sc_hd__o21ai_1 _22445_ (.A1(_06205_),
    .A2(_06233_),
    .B1(net1633),
    .Y(_01584_));
 sky130_fd_sc_hd__a211o_1 _22446_ (.A1(_05564_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06199_),
    .X(_06235_));
 sky130_fd_sc_hd__nand2_1 _22447_ (.A(_06177_),
    .B(net622),
    .Y(_06236_));
 sky130_fd_sc_hd__o21ai_1 _22448_ (.A1(_06205_),
    .A2(_06235_),
    .B1(net623),
    .Y(_01585_));
 sky130_fd_sc_hd__a211o_1 _22449_ (.A1(_05567_),
    .A2(_06179_),
    .B1(_06210_),
    .C1(_06202_),
    .X(_06237_));
 sky130_fd_sc_hd__nand2_1 _22450_ (.A(_06177_),
    .B(net660),
    .Y(_06238_));
 sky130_fd_sc_hd__o21ai_1 _22451_ (.A1(_06205_),
    .A2(_06237_),
    .B1(net661),
    .Y(_01586_));
 sky130_fd_sc_hd__and3_4 _22452_ (.A(_12173_),
    .B(\line_cache_idx[7] ),
    .C(_12303_),
    .X(_06239_));
 sky130_fd_sc_hd__nand2_1 _22453_ (.A(_06239_),
    .B(_04104_),
    .Y(_06240_));
 sky130_fd_sc_hd__a21bo_1 _22454_ (.A1(_06240_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_8 _22455_ (.A(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__mux2_1 _22456_ (.A0(_05318_),
    .A1(net3448),
    .S(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _22457_ (.A(_06243_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _22458_ (.A0(_05324_),
    .A1(net2987),
    .S(_06242_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _22459_ (.A(_06244_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _22460_ (.A0(_05326_),
    .A1(net3656),
    .S(_06242_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _22461_ (.A(_06245_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _22462_ (.A0(_05328_),
    .A1(net3288),
    .S(_06242_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _22463_ (.A(_06246_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _22464_ (.A0(_05330_),
    .A1(net3234),
    .S(_06242_),
    .X(_06247_));
 sky130_fd_sc_hd__clkbuf_1 _22465_ (.A(_06247_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _22466_ (.A0(_05332_),
    .A1(net2602),
    .S(_06242_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _22467_ (.A(_06248_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _22468_ (.A0(_05334_),
    .A1(net2397),
    .S(_06242_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _22469_ (.A(_06249_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _22470_ (.A0(_05336_),
    .A1(net3223),
    .S(_06242_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _22471_ (.A(_06250_),
    .X(_01594_));
 sky130_fd_sc_hd__buf_4 _22472_ (.A(_06240_),
    .X(_06251_));
 sky130_fd_sc_hd__buf_4 _22473_ (.A(_05183_),
    .X(_06252_));
 sky130_fd_sc_hd__buf_4 _22474_ (.A(_06240_),
    .X(_06253_));
 sky130_fd_sc_hd__nand2_1 _22475_ (.A(_06253_),
    .B(_05010_),
    .Y(_06254_));
 sky130_fd_sc_hd__o211a_1 _22476_ (.A1(_05095_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__mux2_1 _22477_ (.A0(_06255_),
    .A1(net3299),
    .S(_06242_),
    .X(_06256_));
 sky130_fd_sc_hd__clkbuf_1 _22478_ (.A(_06256_),
    .X(_01595_));
 sky130_fd_sc_hd__nand2_1 _22479_ (.A(_06253_),
    .B(_05014_),
    .Y(_06257_));
 sky130_fd_sc_hd__o211a_1 _22480_ (.A1(_05101_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__mux2_1 _22481_ (.A0(_06258_),
    .A1(net2458),
    .S(_06242_),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _22482_ (.A(_06259_),
    .X(_01596_));
 sky130_fd_sc_hd__nand2_1 _22483_ (.A(_06253_),
    .B(_05018_),
    .Y(_06260_));
 sky130_fd_sc_hd__o211a_1 _22484_ (.A1(_05105_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__mux2_1 _22485_ (.A0(_06261_),
    .A1(net2443),
    .S(_06242_),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _22486_ (.A(_06262_),
    .X(_01597_));
 sky130_fd_sc_hd__nand2_1 _22487_ (.A(_06253_),
    .B(_05022_),
    .Y(_06263_));
 sky130_fd_sc_hd__o211a_1 _22488_ (.A1(_05109_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__mux2_1 _22489_ (.A0(_06264_),
    .A1(net2648),
    .S(_06242_),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_1 _22490_ (.A(_06265_),
    .X(_01598_));
 sky130_fd_sc_hd__nand2_1 _22491_ (.A(_06253_),
    .B(_05026_),
    .Y(_06266_));
 sky130_fd_sc_hd__o211a_1 _22492_ (.A1(_05113_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__mux2_1 _22493_ (.A0(_06267_),
    .A1(net2801),
    .S(_06242_),
    .X(_06268_));
 sky130_fd_sc_hd__clkbuf_1 _22494_ (.A(_06268_),
    .X(_01599_));
 sky130_fd_sc_hd__nand2_1 _22495_ (.A(_06253_),
    .B(_05030_),
    .Y(_06269_));
 sky130_fd_sc_hd__o211a_1 _22496_ (.A1(_05117_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__mux2_1 _22497_ (.A0(_06270_),
    .A1(net2466),
    .S(_06242_),
    .X(_06271_));
 sky130_fd_sc_hd__clkbuf_1 _22498_ (.A(_06271_),
    .X(_01600_));
 sky130_fd_sc_hd__nand2_1 _22499_ (.A(_06253_),
    .B(_05034_),
    .Y(_06272_));
 sky130_fd_sc_hd__o211a_1 _22500_ (.A1(_05121_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__mux2_1 _22501_ (.A0(_06273_),
    .A1(net3081),
    .S(_06242_),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_1 _22502_ (.A(_06274_),
    .X(_01601_));
 sky130_fd_sc_hd__nand2_1 _22503_ (.A(_06253_),
    .B(_05038_),
    .Y(_06275_));
 sky130_fd_sc_hd__o211a_1 _22504_ (.A1(_05125_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__mux2_1 _22505_ (.A0(_06276_),
    .A1(net3043),
    .S(_06242_),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_1 _22506_ (.A(_06277_),
    .X(_01602_));
 sky130_fd_sc_hd__o211a_1 _22507_ (.A1(_05129_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06254_),
    .X(_06278_));
 sky130_fd_sc_hd__clkbuf_8 _22508_ (.A(_06241_),
    .X(_06279_));
 sky130_fd_sc_hd__mux2_1 _22509_ (.A0(_06278_),
    .A1(net2992),
    .S(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__clkbuf_1 _22510_ (.A(_06280_),
    .X(_01603_));
 sky130_fd_sc_hd__o211a_1 _22511_ (.A1(_05134_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06257_),
    .X(_06281_));
 sky130_fd_sc_hd__mux2_1 _22512_ (.A0(_06281_),
    .A1(net3635),
    .S(_06279_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _22513_ (.A(_06282_),
    .X(_01604_));
 sky130_fd_sc_hd__o211a_1 _22514_ (.A1(_05137_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06260_),
    .X(_06283_));
 sky130_fd_sc_hd__mux2_1 _22515_ (.A0(_06283_),
    .A1(net3743),
    .S(_06279_),
    .X(_06284_));
 sky130_fd_sc_hd__clkbuf_1 _22516_ (.A(_06284_),
    .X(_01605_));
 sky130_fd_sc_hd__o211a_1 _22517_ (.A1(_05140_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06263_),
    .X(_06285_));
 sky130_fd_sc_hd__mux2_1 _22518_ (.A0(_06285_),
    .A1(net2673),
    .S(_06279_),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _22519_ (.A(_06286_),
    .X(_01606_));
 sky130_fd_sc_hd__o211a_1 _22520_ (.A1(_05143_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06266_),
    .X(_06287_));
 sky130_fd_sc_hd__mux2_1 _22521_ (.A0(_06287_),
    .A1(net3754),
    .S(_06279_),
    .X(_06288_));
 sky130_fd_sc_hd__clkbuf_1 _22522_ (.A(_06288_),
    .X(_01607_));
 sky130_fd_sc_hd__o211a_1 _22523_ (.A1(_05146_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06269_),
    .X(_06289_));
 sky130_fd_sc_hd__mux2_1 _22524_ (.A0(_06289_),
    .A1(net3722),
    .S(_06279_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _22525_ (.A(_06290_),
    .X(_01608_));
 sky130_fd_sc_hd__o211a_1 _22526_ (.A1(_05149_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06272_),
    .X(_06291_));
 sky130_fd_sc_hd__mux2_1 _22527_ (.A0(_06291_),
    .A1(net3686),
    .S(_06279_),
    .X(_06292_));
 sky130_fd_sc_hd__clkbuf_1 _22528_ (.A(_06292_),
    .X(_01609_));
 sky130_fd_sc_hd__o211a_1 _22529_ (.A1(_05152_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06275_),
    .X(_06293_));
 sky130_fd_sc_hd__mux2_1 _22530_ (.A0(_06293_),
    .A1(net3009),
    .S(_06279_),
    .X(_06294_));
 sky130_fd_sc_hd__clkbuf_1 _22531_ (.A(_06294_),
    .X(_01610_));
 sky130_fd_sc_hd__clkbuf_8 _22532_ (.A(_05183_),
    .X(_06295_));
 sky130_fd_sc_hd__o211a_1 _22533_ (.A1(_05059_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06254_),
    .X(_06296_));
 sky130_fd_sc_hd__mux2_1 _22534_ (.A0(_06296_),
    .A1(net2196),
    .S(_06279_),
    .X(_06297_));
 sky130_fd_sc_hd__clkbuf_1 _22535_ (.A(_06297_),
    .X(_01611_));
 sky130_fd_sc_hd__o211a_1 _22536_ (.A1(_05063_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06257_),
    .X(_06298_));
 sky130_fd_sc_hd__mux2_1 _22537_ (.A0(_06298_),
    .A1(net3723),
    .S(_06279_),
    .X(_06299_));
 sky130_fd_sc_hd__clkbuf_1 _22538_ (.A(_06299_),
    .X(_01612_));
 sky130_fd_sc_hd__o211a_1 _22539_ (.A1(_05066_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06260_),
    .X(_06300_));
 sky130_fd_sc_hd__mux2_1 _22540_ (.A0(_06300_),
    .A1(net3672),
    .S(_06279_),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_1 _22541_ (.A(_06301_),
    .X(_01613_));
 sky130_fd_sc_hd__o211a_1 _22542_ (.A1(_05069_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06263_),
    .X(_06302_));
 sky130_fd_sc_hd__mux2_1 _22543_ (.A0(_06302_),
    .A1(net2913),
    .S(_06279_),
    .X(_06303_));
 sky130_fd_sc_hd__clkbuf_1 _22544_ (.A(_06303_),
    .X(_01614_));
 sky130_fd_sc_hd__o211a_1 _22545_ (.A1(_05072_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06266_),
    .X(_06304_));
 sky130_fd_sc_hd__mux2_1 _22546_ (.A0(_06304_),
    .A1(net3633),
    .S(_06279_),
    .X(_06305_));
 sky130_fd_sc_hd__clkbuf_1 _22547_ (.A(_06305_),
    .X(_01615_));
 sky130_fd_sc_hd__o211a_1 _22548_ (.A1(_05075_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06269_),
    .X(_06306_));
 sky130_fd_sc_hd__mux2_1 _22549_ (.A0(_06306_),
    .A1(net3733),
    .S(_06279_),
    .X(_06307_));
 sky130_fd_sc_hd__clkbuf_1 _22550_ (.A(_06307_),
    .X(_01616_));
 sky130_fd_sc_hd__o211a_1 _22551_ (.A1(_05078_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06272_),
    .X(_06308_));
 sky130_fd_sc_hd__mux2_1 _22552_ (.A0(_06308_),
    .A1(net3663),
    .S(_06279_),
    .X(_06309_));
 sky130_fd_sc_hd__clkbuf_1 _22553_ (.A(_06309_),
    .X(_01617_));
 sky130_fd_sc_hd__o211a_1 _22554_ (.A1(_05081_),
    .A2(_06253_),
    .B1(_06295_),
    .C1(_06275_),
    .X(_06310_));
 sky130_fd_sc_hd__mux2_1 _22555_ (.A0(_06310_),
    .A1(net3178),
    .S(_06279_),
    .X(_06311_));
 sky130_fd_sc_hd__clkbuf_1 _22556_ (.A(_06311_),
    .X(_01618_));
 sky130_fd_sc_hd__nand2_1 _22557_ (.A(_06239_),
    .B(_04183_),
    .Y(_06312_));
 sky130_fd_sc_hd__a21bo_1 _22558_ (.A1(_06312_),
    .A2(_03813_),
    .B1_N(_03739_),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_8 _22559_ (.A(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_1 _22560_ (.A0(_05318_),
    .A1(net2259),
    .S(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _22561_ (.A(_06315_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _22562_ (.A0(_05324_),
    .A1(net2268),
    .S(_06314_),
    .X(_06316_));
 sky130_fd_sc_hd__clkbuf_1 _22563_ (.A(_06316_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _22564_ (.A0(_05326_),
    .A1(net2659),
    .S(_06314_),
    .X(_06317_));
 sky130_fd_sc_hd__clkbuf_1 _22565_ (.A(_06317_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _22566_ (.A0(_05328_),
    .A1(net2331),
    .S(_06314_),
    .X(_06318_));
 sky130_fd_sc_hd__clkbuf_1 _22567_ (.A(_06318_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _22568_ (.A0(_05330_),
    .A1(net2969),
    .S(_06314_),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_1 _22569_ (.A(_06319_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _22570_ (.A0(_05332_),
    .A1(net2784),
    .S(_06314_),
    .X(_06320_));
 sky130_fd_sc_hd__clkbuf_1 _22571_ (.A(_06320_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _22572_ (.A0(_05334_),
    .A1(net3137),
    .S(_06314_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _22573_ (.A(_06321_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _22574_ (.A0(_05336_),
    .A1(net2252),
    .S(_06314_),
    .X(_06322_));
 sky130_fd_sc_hd__clkbuf_1 _22575_ (.A(_06322_),
    .X(_01626_));
 sky130_fd_sc_hd__buf_4 _22576_ (.A(_06312_),
    .X(_06323_));
 sky130_fd_sc_hd__buf_4 _22577_ (.A(_06312_),
    .X(_06324_));
 sky130_fd_sc_hd__nand2_1 _22578_ (.A(_06324_),
    .B(_05010_),
    .Y(_06325_));
 sky130_fd_sc_hd__o211a_1 _22579_ (.A1(_05095_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__mux2_1 _22580_ (.A0(_06326_),
    .A1(net2024),
    .S(_06314_),
    .X(_06327_));
 sky130_fd_sc_hd__clkbuf_1 _22581_ (.A(_06327_),
    .X(_01627_));
 sky130_fd_sc_hd__nand2_1 _22582_ (.A(_06324_),
    .B(_05014_),
    .Y(_06328_));
 sky130_fd_sc_hd__o211a_1 _22583_ (.A1(_05101_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__mux2_1 _22584_ (.A0(_06329_),
    .A1(net2139),
    .S(_06314_),
    .X(_06330_));
 sky130_fd_sc_hd__clkbuf_1 _22585_ (.A(_06330_),
    .X(_01628_));
 sky130_fd_sc_hd__nand2_1 _22586_ (.A(_06324_),
    .B(_05018_),
    .Y(_06331_));
 sky130_fd_sc_hd__o211a_1 _22587_ (.A1(_05105_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__mux2_1 _22588_ (.A0(_06332_),
    .A1(net2236),
    .S(_06314_),
    .X(_06333_));
 sky130_fd_sc_hd__clkbuf_1 _22589_ (.A(_06333_),
    .X(_01629_));
 sky130_fd_sc_hd__nand2_1 _22590_ (.A(_06324_),
    .B(_05022_),
    .Y(_06334_));
 sky130_fd_sc_hd__o211a_1 _22591_ (.A1(_05109_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__mux2_1 _22592_ (.A0(_06335_),
    .A1(net2282),
    .S(_06314_),
    .X(_06336_));
 sky130_fd_sc_hd__clkbuf_1 _22593_ (.A(_06336_),
    .X(_01630_));
 sky130_fd_sc_hd__nand2_1 _22594_ (.A(_06324_),
    .B(_05026_),
    .Y(_06337_));
 sky130_fd_sc_hd__o211a_1 _22595_ (.A1(_05113_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__mux2_1 _22596_ (.A0(_06338_),
    .A1(net2155),
    .S(_06314_),
    .X(_06339_));
 sky130_fd_sc_hd__clkbuf_1 _22597_ (.A(_06339_),
    .X(_01631_));
 sky130_fd_sc_hd__nand2_1 _22598_ (.A(_06324_),
    .B(_05030_),
    .Y(_06340_));
 sky130_fd_sc_hd__o211a_1 _22599_ (.A1(_05117_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__mux2_1 _22600_ (.A0(_06341_),
    .A1(net2074),
    .S(_06314_),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_1 _22601_ (.A(_06342_),
    .X(_01632_));
 sky130_fd_sc_hd__nand2_1 _22602_ (.A(_06324_),
    .B(_05034_),
    .Y(_06343_));
 sky130_fd_sc_hd__o211a_1 _22603_ (.A1(_05121_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__mux2_1 _22604_ (.A0(_06344_),
    .A1(net2084),
    .S(_06314_),
    .X(_06345_));
 sky130_fd_sc_hd__clkbuf_1 _22605_ (.A(_06345_),
    .X(_01633_));
 sky130_fd_sc_hd__nand2_1 _22606_ (.A(_06324_),
    .B(_05038_),
    .Y(_06346_));
 sky130_fd_sc_hd__o211a_1 _22607_ (.A1(_05125_),
    .A2(_06323_),
    .B1(_06295_),
    .C1(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__mux2_1 _22608_ (.A0(_06347_),
    .A1(net2098),
    .S(_06314_),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_1 _22609_ (.A(_06348_),
    .X(_01634_));
 sky130_fd_sc_hd__buf_4 _22610_ (.A(_05183_),
    .X(_06349_));
 sky130_fd_sc_hd__o211a_1 _22611_ (.A1(_05129_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06325_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_8 _22612_ (.A(_06313_),
    .X(_06351_));
 sky130_fd_sc_hd__mux2_1 _22613_ (.A0(_06350_),
    .A1(net2564),
    .S(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__clkbuf_1 _22614_ (.A(_06352_),
    .X(_01635_));
 sky130_fd_sc_hd__o211a_1 _22615_ (.A1(_05134_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06328_),
    .X(_06353_));
 sky130_fd_sc_hd__mux2_1 _22616_ (.A0(_06353_),
    .A1(net2108),
    .S(_06351_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _22617_ (.A(_06354_),
    .X(_01636_));
 sky130_fd_sc_hd__o211a_1 _22618_ (.A1(_05137_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06331_),
    .X(_06355_));
 sky130_fd_sc_hd__mux2_1 _22619_ (.A0(_06355_),
    .A1(net2078),
    .S(_06351_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _22620_ (.A(_06356_),
    .X(_01637_));
 sky130_fd_sc_hd__o211a_1 _22621_ (.A1(_05140_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06334_),
    .X(_06357_));
 sky130_fd_sc_hd__mux2_1 _22622_ (.A0(_06357_),
    .A1(net2257),
    .S(_06351_),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_1 _22623_ (.A(_06358_),
    .X(_01638_));
 sky130_fd_sc_hd__o211a_1 _22624_ (.A1(_05143_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06337_),
    .X(_06359_));
 sky130_fd_sc_hd__mux2_1 _22625_ (.A0(_06359_),
    .A1(net2064),
    .S(_06351_),
    .X(_06360_));
 sky130_fd_sc_hd__clkbuf_1 _22626_ (.A(_06360_),
    .X(_01639_));
 sky130_fd_sc_hd__o211a_1 _22627_ (.A1(_05146_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06340_),
    .X(_06361_));
 sky130_fd_sc_hd__mux2_1 _22628_ (.A0(_06361_),
    .A1(net2068),
    .S(_06351_),
    .X(_06362_));
 sky130_fd_sc_hd__clkbuf_1 _22629_ (.A(_06362_),
    .X(_01640_));
 sky130_fd_sc_hd__o211a_1 _22630_ (.A1(_05149_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06343_),
    .X(_06363_));
 sky130_fd_sc_hd__mux2_1 _22631_ (.A0(_06363_),
    .A1(net2082),
    .S(_06351_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_1 _22632_ (.A(_06364_),
    .X(_01641_));
 sky130_fd_sc_hd__o211a_1 _22633_ (.A1(_05152_),
    .A2(_06323_),
    .B1(_06349_),
    .C1(_06346_),
    .X(_06365_));
 sky130_fd_sc_hd__mux2_1 _22634_ (.A0(_06365_),
    .A1(net2131),
    .S(_06351_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _22635_ (.A(_06366_),
    .X(_01642_));
 sky130_fd_sc_hd__o211a_1 _22636_ (.A1(_05059_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06325_),
    .X(_06367_));
 sky130_fd_sc_hd__mux2_1 _22637_ (.A0(_06367_),
    .A1(net2035),
    .S(_06351_),
    .X(_06368_));
 sky130_fd_sc_hd__clkbuf_1 _22638_ (.A(_06368_),
    .X(_01643_));
 sky130_fd_sc_hd__o211a_1 _22639_ (.A1(_05063_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06328_),
    .X(_06369_));
 sky130_fd_sc_hd__mux2_1 _22640_ (.A0(_06369_),
    .A1(net2177),
    .S(_06351_),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_1 _22641_ (.A(_06370_),
    .X(_01644_));
 sky130_fd_sc_hd__o211a_1 _22642_ (.A1(_05066_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06331_),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_1 _22643_ (.A0(_06371_),
    .A1(net3674),
    .S(_06351_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _22644_ (.A(_06372_),
    .X(_01645_));
 sky130_fd_sc_hd__o211a_1 _22645_ (.A1(_05069_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06334_),
    .X(_06373_));
 sky130_fd_sc_hd__mux2_1 _22646_ (.A0(_06373_),
    .A1(net3616),
    .S(_06351_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_1 _22647_ (.A(_06374_),
    .X(_01646_));
 sky130_fd_sc_hd__o211a_1 _22648_ (.A1(_05072_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06337_),
    .X(_06375_));
 sky130_fd_sc_hd__mux2_1 _22649_ (.A0(_06375_),
    .A1(net2714),
    .S(_06351_),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_1 _22650_ (.A(_06376_),
    .X(_01647_));
 sky130_fd_sc_hd__o211a_1 _22651_ (.A1(_05075_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06340_),
    .X(_06377_));
 sky130_fd_sc_hd__mux2_1 _22652_ (.A0(_06377_),
    .A1(net3657),
    .S(_06351_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _22653_ (.A(_06378_),
    .X(_01648_));
 sky130_fd_sc_hd__o211a_1 _22654_ (.A1(_05078_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06343_),
    .X(_06379_));
 sky130_fd_sc_hd__mux2_1 _22655_ (.A0(_06379_),
    .A1(net3587),
    .S(_06351_),
    .X(_06380_));
 sky130_fd_sc_hd__clkbuf_1 _22656_ (.A(_06380_),
    .X(_01649_));
 sky130_fd_sc_hd__o211a_1 _22657_ (.A1(_05081_),
    .A2(_06324_),
    .B1(_06349_),
    .C1(_06346_),
    .X(_06381_));
 sky130_fd_sc_hd__mux2_1 _22658_ (.A0(_06381_),
    .A1(net3602),
    .S(_06351_),
    .X(_06382_));
 sky130_fd_sc_hd__clkbuf_1 _22659_ (.A(_06382_),
    .X(_01650_));
 sky130_fd_sc_hd__nand2_1 _22660_ (.A(_06239_),
    .B(_04257_),
    .Y(_06383_));
 sky130_fd_sc_hd__buf_6 _22661_ (.A(_12189_),
    .X(_06384_));
 sky130_fd_sc_hd__a21bo_1 _22662_ (.A1(_06383_),
    .A2(_03813_),
    .B1_N(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_8 _22663_ (.A(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__mux2_1 _22664_ (.A0(_05318_),
    .A1(net2523),
    .S(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__clkbuf_1 _22665_ (.A(_06387_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _22666_ (.A0(_05324_),
    .A1(net3726),
    .S(_06386_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_1 _22667_ (.A(_06388_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _22668_ (.A0(_05326_),
    .A1(net2510),
    .S(_06386_),
    .X(_06389_));
 sky130_fd_sc_hd__clkbuf_1 _22669_ (.A(_06389_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _22670_ (.A0(_05328_),
    .A1(net3109),
    .S(_06386_),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_1 _22671_ (.A(_06390_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _22672_ (.A0(_05330_),
    .A1(net3031),
    .S(_06386_),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_1 _22673_ (.A(_06391_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _22674_ (.A0(_05332_),
    .A1(net3513),
    .S(_06386_),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _22675_ (.A(_06392_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _22676_ (.A0(_05334_),
    .A1(net3770),
    .S(_06386_),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _22677_ (.A(_06393_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _22678_ (.A0(_05336_),
    .A1(net3308),
    .S(_06386_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _22679_ (.A(_06394_),
    .X(_01658_));
 sky130_fd_sc_hd__buf_4 _22680_ (.A(_06383_),
    .X(_06395_));
 sky130_fd_sc_hd__buf_4 _22681_ (.A(_05183_),
    .X(_06396_));
 sky130_fd_sc_hd__buf_4 _22682_ (.A(_06383_),
    .X(_06397_));
 sky130_fd_sc_hd__nand2_1 _22683_ (.A(_06397_),
    .B(_05010_),
    .Y(_06398_));
 sky130_fd_sc_hd__o211a_1 _22684_ (.A1(_05095_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__mux2_1 _22685_ (.A0(_06399_),
    .A1(net2465),
    .S(_06386_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_1 _22686_ (.A(_06400_),
    .X(_01659_));
 sky130_fd_sc_hd__nand2_1 _22687_ (.A(_06397_),
    .B(_05014_),
    .Y(_06401_));
 sky130_fd_sc_hd__o211a_1 _22688_ (.A1(_05101_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__mux2_1 _22689_ (.A0(_06402_),
    .A1(net2839),
    .S(_06386_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _22690_ (.A(_06403_),
    .X(_01660_));
 sky130_fd_sc_hd__nand2_1 _22691_ (.A(_06397_),
    .B(_05018_),
    .Y(_06404_));
 sky130_fd_sc_hd__o211a_1 _22692_ (.A1(_05105_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__mux2_1 _22693_ (.A0(_06405_),
    .A1(net2288),
    .S(_06386_),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_1 _22694_ (.A(_06406_),
    .X(_01661_));
 sky130_fd_sc_hd__nand2_1 _22695_ (.A(_06397_),
    .B(_05022_),
    .Y(_06407_));
 sky130_fd_sc_hd__o211a_1 _22696_ (.A1(_05109_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__mux2_1 _22697_ (.A0(_06408_),
    .A1(net2292),
    .S(_06386_),
    .X(_06409_));
 sky130_fd_sc_hd__clkbuf_1 _22698_ (.A(_06409_),
    .X(_01662_));
 sky130_fd_sc_hd__nand2_1 _22699_ (.A(_06397_),
    .B(_05026_),
    .Y(_06410_));
 sky130_fd_sc_hd__o211a_1 _22700_ (.A1(_05113_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__mux2_1 _22701_ (.A0(_06411_),
    .A1(net3244),
    .S(_06386_),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_1 _22702_ (.A(_06412_),
    .X(_01663_));
 sky130_fd_sc_hd__nand2_1 _22703_ (.A(_06397_),
    .B(_05030_),
    .Y(_06413_));
 sky130_fd_sc_hd__o211a_1 _22704_ (.A1(_05117_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__mux2_1 _22705_ (.A0(_06414_),
    .A1(net3263),
    .S(_06386_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _22706_ (.A(_06415_),
    .X(_01664_));
 sky130_fd_sc_hd__nand2_1 _22707_ (.A(_06397_),
    .B(_05034_),
    .Y(_06416_));
 sky130_fd_sc_hd__o211a_1 _22708_ (.A1(_05121_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__mux2_1 _22709_ (.A0(_06417_),
    .A1(net2653),
    .S(_06386_),
    .X(_06418_));
 sky130_fd_sc_hd__clkbuf_1 _22710_ (.A(_06418_),
    .X(_01665_));
 sky130_fd_sc_hd__nand2_1 _22711_ (.A(_06397_),
    .B(_05038_),
    .Y(_06419_));
 sky130_fd_sc_hd__o211a_1 _22712_ (.A1(_05125_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__mux2_1 _22713_ (.A0(_06420_),
    .A1(net2721),
    .S(_06386_),
    .X(_06421_));
 sky130_fd_sc_hd__clkbuf_1 _22714_ (.A(_06421_),
    .X(_01666_));
 sky130_fd_sc_hd__o211a_1 _22715_ (.A1(_05129_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06398_),
    .X(_06422_));
 sky130_fd_sc_hd__clkbuf_8 _22716_ (.A(_06385_),
    .X(_06423_));
 sky130_fd_sc_hd__mux2_1 _22717_ (.A0(_06422_),
    .A1(net3869),
    .S(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__clkbuf_1 _22718_ (.A(_06424_),
    .X(_01667_));
 sky130_fd_sc_hd__o211a_1 _22719_ (.A1(_05134_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06401_),
    .X(_06425_));
 sky130_fd_sc_hd__mux2_1 _22720_ (.A0(_06425_),
    .A1(net2392),
    .S(_06423_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _22721_ (.A(_06426_),
    .X(_01668_));
 sky130_fd_sc_hd__o211a_1 _22722_ (.A1(_05137_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06404_),
    .X(_06427_));
 sky130_fd_sc_hd__mux2_1 _22723_ (.A0(_06427_),
    .A1(net3147),
    .S(_06423_),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_1 _22724_ (.A(_06428_),
    .X(_01669_));
 sky130_fd_sc_hd__o211a_1 _22725_ (.A1(_05140_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06407_),
    .X(_06429_));
 sky130_fd_sc_hd__mux2_1 _22726_ (.A0(_06429_),
    .A1(net2705),
    .S(_06423_),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_1 _22727_ (.A(_06430_),
    .X(_01670_));
 sky130_fd_sc_hd__o211a_1 _22728_ (.A1(_05143_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06410_),
    .X(_06431_));
 sky130_fd_sc_hd__mux2_1 _22729_ (.A0(_06431_),
    .A1(net2822),
    .S(_06423_),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_1 _22730_ (.A(_06432_),
    .X(_01671_));
 sky130_fd_sc_hd__o211a_1 _22731_ (.A1(_05146_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06413_),
    .X(_06433_));
 sky130_fd_sc_hd__mux2_1 _22732_ (.A0(_06433_),
    .A1(net2574),
    .S(_06423_),
    .X(_06434_));
 sky130_fd_sc_hd__clkbuf_1 _22733_ (.A(_06434_),
    .X(_01672_));
 sky130_fd_sc_hd__o211a_1 _22734_ (.A1(_05149_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06416_),
    .X(_06435_));
 sky130_fd_sc_hd__mux2_1 _22735_ (.A0(_06435_),
    .A1(net3626),
    .S(_06423_),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_1 _22736_ (.A(_06436_),
    .X(_01673_));
 sky130_fd_sc_hd__o211a_1 _22737_ (.A1(_05152_),
    .A2(_06395_),
    .B1(_06396_),
    .C1(_06419_),
    .X(_06437_));
 sky130_fd_sc_hd__mux2_1 _22738_ (.A0(_06437_),
    .A1(net3642),
    .S(_06423_),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_1 _22739_ (.A(_06438_),
    .X(_01674_));
 sky130_fd_sc_hd__clkbuf_8 _22740_ (.A(_05183_),
    .X(_06439_));
 sky130_fd_sc_hd__o211a_1 _22741_ (.A1(_05059_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06398_),
    .X(_06440_));
 sky130_fd_sc_hd__mux2_1 _22742_ (.A0(_06440_),
    .A1(net3898),
    .S(_06423_),
    .X(_06441_));
 sky130_fd_sc_hd__clkbuf_1 _22743_ (.A(_06441_),
    .X(_01675_));
 sky130_fd_sc_hd__o211a_1 _22744_ (.A1(_05063_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06401_),
    .X(_06442_));
 sky130_fd_sc_hd__mux2_1 _22745_ (.A0(_06442_),
    .A1(net3321),
    .S(_06423_),
    .X(_06443_));
 sky130_fd_sc_hd__clkbuf_1 _22746_ (.A(_06443_),
    .X(_01676_));
 sky130_fd_sc_hd__o211a_1 _22747_ (.A1(_05066_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06404_),
    .X(_06444_));
 sky130_fd_sc_hd__mux2_1 _22748_ (.A0(_06444_),
    .A1(net2537),
    .S(_06423_),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_1 _22749_ (.A(_06445_),
    .X(_01677_));
 sky130_fd_sc_hd__o211a_1 _22750_ (.A1(_05069_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06407_),
    .X(_06446_));
 sky130_fd_sc_hd__mux2_1 _22751_ (.A0(_06446_),
    .A1(net2732),
    .S(_06423_),
    .X(_06447_));
 sky130_fd_sc_hd__clkbuf_1 _22752_ (.A(_06447_),
    .X(_01678_));
 sky130_fd_sc_hd__o211a_1 _22753_ (.A1(_05072_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06410_),
    .X(_06448_));
 sky130_fd_sc_hd__mux2_1 _22754_ (.A0(_06448_),
    .A1(net2427),
    .S(_06423_),
    .X(_06449_));
 sky130_fd_sc_hd__clkbuf_1 _22755_ (.A(_06449_),
    .X(_01679_));
 sky130_fd_sc_hd__o211a_1 _22756_ (.A1(_05075_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06413_),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_1 _22757_ (.A0(_06450_),
    .A1(net3158),
    .S(_06423_),
    .X(_06451_));
 sky130_fd_sc_hd__clkbuf_1 _22758_ (.A(_06451_),
    .X(_01680_));
 sky130_fd_sc_hd__o211a_1 _22759_ (.A1(_05078_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06416_),
    .X(_06452_));
 sky130_fd_sc_hd__mux2_1 _22760_ (.A0(_06452_),
    .A1(net3670),
    .S(_06423_),
    .X(_06453_));
 sky130_fd_sc_hd__clkbuf_1 _22761_ (.A(_06453_),
    .X(_01681_));
 sky130_fd_sc_hd__o211a_1 _22762_ (.A1(_05081_),
    .A2(_06397_),
    .B1(_06439_),
    .C1(_06419_),
    .X(_06454_));
 sky130_fd_sc_hd__mux2_1 _22763_ (.A0(_06454_),
    .A1(net3702),
    .S(_06423_),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_1 _22764_ (.A(_06455_),
    .X(_01682_));
 sky130_fd_sc_hd__nand2_1 _22765_ (.A(_06239_),
    .B(_04333_),
    .Y(_06456_));
 sky130_fd_sc_hd__inv_2 _22766_ (.A(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__o21ai_4 _22767_ (.A1(_05471_),
    .A2(_06457_),
    .B1(_06020_),
    .Y(_06458_));
 sky130_fd_sc_hd__mux2_1 _22768_ (.A0(_05318_),
    .A1(net2353),
    .S(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__clkbuf_1 _22769_ (.A(_06459_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _22770_ (.A0(_05324_),
    .A1(net3584),
    .S(_06458_),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_1 _22771_ (.A(_06460_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _22772_ (.A0(_05326_),
    .A1(net2840),
    .S(_06458_),
    .X(_06461_));
 sky130_fd_sc_hd__clkbuf_1 _22773_ (.A(_06461_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _22774_ (.A0(_05328_),
    .A1(net2586),
    .S(_06458_),
    .X(_06462_));
 sky130_fd_sc_hd__clkbuf_1 _22775_ (.A(_06462_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _22776_ (.A0(_05330_),
    .A1(net3554),
    .S(_06458_),
    .X(_06463_));
 sky130_fd_sc_hd__clkbuf_1 _22777_ (.A(_06463_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _22778_ (.A0(_05332_),
    .A1(net3509),
    .S(_06458_),
    .X(_06464_));
 sky130_fd_sc_hd__clkbuf_1 _22779_ (.A(_06464_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _22780_ (.A0(_05334_),
    .A1(net2582),
    .S(_06458_),
    .X(_06465_));
 sky130_fd_sc_hd__clkbuf_1 _22781_ (.A(_06465_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _22782_ (.A0(_05336_),
    .A1(net2629),
    .S(_06458_),
    .X(_06466_));
 sky130_fd_sc_hd__clkbuf_1 _22783_ (.A(_06466_),
    .X(_01690_));
 sky130_fd_sc_hd__buf_4 _22784_ (.A(_06458_),
    .X(_06467_));
 sky130_fd_sc_hd__buf_4 _22785_ (.A(_06457_),
    .X(_06468_));
 sky130_fd_sc_hd__buf_4 _22786_ (.A(_06457_),
    .X(_06469_));
 sky130_fd_sc_hd__nor2_1 _22787_ (.A(_05583_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__a211o_1 _22788_ (.A1(_05484_),
    .A2(_06468_),
    .B1(_06210_),
    .C1(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__buf_4 _22789_ (.A(_06458_),
    .X(_06472_));
 sky130_fd_sc_hd__nand2_1 _22790_ (.A(_06472_),
    .B(net1412),
    .Y(_06473_));
 sky130_fd_sc_hd__o21ai_1 _22791_ (.A1(_06467_),
    .A2(_06471_),
    .B1(net1413),
    .Y(_01691_));
 sky130_fd_sc_hd__nor2_1 _22792_ (.A(_05589_),
    .B(_06469_),
    .Y(_06474_));
 sky130_fd_sc_hd__a211o_1 _22793_ (.A1(_05491_),
    .A2(_06468_),
    .B1(_06210_),
    .C1(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__nand2_1 _22794_ (.A(_06472_),
    .B(net1510),
    .Y(_06476_));
 sky130_fd_sc_hd__o21ai_1 _22795_ (.A1(_06467_),
    .A2(_06475_),
    .B1(net1511),
    .Y(_01692_));
 sky130_fd_sc_hd__buf_4 _22796_ (.A(_05892_),
    .X(_06477_));
 sky130_fd_sc_hd__nor2_1 _22797_ (.A(_05593_),
    .B(_06469_),
    .Y(_06478_));
 sky130_fd_sc_hd__a211o_1 _22798_ (.A1(_05495_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__nand2_1 _22799_ (.A(_06472_),
    .B(net1168),
    .Y(_06480_));
 sky130_fd_sc_hd__o21ai_1 _22800_ (.A1(_06467_),
    .A2(_06479_),
    .B1(net1169),
    .Y(_01693_));
 sky130_fd_sc_hd__nor2_1 _22801_ (.A(_05597_),
    .B(_06469_),
    .Y(_06481_));
 sky130_fd_sc_hd__a211o_1 _22802_ (.A1(_05500_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__nand2_1 _22803_ (.A(_06472_),
    .B(net1654),
    .Y(_06483_));
 sky130_fd_sc_hd__o21ai_1 _22804_ (.A1(_06467_),
    .A2(_06482_),
    .B1(net1655),
    .Y(_01694_));
 sky130_fd_sc_hd__nor2_1 _22805_ (.A(_05601_),
    .B(_06469_),
    .Y(_06484_));
 sky130_fd_sc_hd__a211o_1 _22806_ (.A1(_05504_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__nand2_1 _22807_ (.A(_06472_),
    .B(net732),
    .Y(_06486_));
 sky130_fd_sc_hd__o21ai_1 _22808_ (.A1(_06467_),
    .A2(_06485_),
    .B1(net733),
    .Y(_01695_));
 sky130_fd_sc_hd__nor2_1 _22809_ (.A(_05605_),
    .B(_06469_),
    .Y(_06487_));
 sky130_fd_sc_hd__a211o_1 _22810_ (.A1(_05508_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06487_),
    .X(_06488_));
 sky130_fd_sc_hd__nand2_1 _22811_ (.A(_06472_),
    .B(net1204),
    .Y(_06489_));
 sky130_fd_sc_hd__o21ai_1 _22812_ (.A1(_06467_),
    .A2(_06488_),
    .B1(net1205),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_1 _22813_ (.A(_05609_),
    .B(_06469_),
    .Y(_06490_));
 sky130_fd_sc_hd__a211o_1 _22814_ (.A1(_05512_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__nand2_1 _22815_ (.A(_06472_),
    .B(net1454),
    .Y(_06492_));
 sky130_fd_sc_hd__o21ai_1 _22816_ (.A1(_06467_),
    .A2(_06491_),
    .B1(net1455),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_1 _22817_ (.A(_05613_),
    .B(_06469_),
    .Y(_06493_));
 sky130_fd_sc_hd__a211o_1 _22818_ (.A1(_05516_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__nand2_1 _22819_ (.A(_06472_),
    .B(net1540),
    .Y(_06495_));
 sky130_fd_sc_hd__o21ai_1 _22820_ (.A1(_06467_),
    .A2(_06494_),
    .B1(net1541),
    .Y(_01698_));
 sky130_fd_sc_hd__buf_4 _22821_ (.A(_06458_),
    .X(_06496_));
 sky130_fd_sc_hd__a211o_1 _22822_ (.A1(_05521_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06470_),
    .X(_06497_));
 sky130_fd_sc_hd__nand2_1 _22823_ (.A(_06472_),
    .B(net634),
    .Y(_06498_));
 sky130_fd_sc_hd__o21ai_1 _22824_ (.A1(_06496_),
    .A2(_06497_),
    .B1(net635),
    .Y(_01699_));
 sky130_fd_sc_hd__a211o_1 _22825_ (.A1(_05524_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06474_),
    .X(_06499_));
 sky130_fd_sc_hd__nand2_1 _22826_ (.A(_06472_),
    .B(net1776),
    .Y(_06500_));
 sky130_fd_sc_hd__o21ai_1 _22827_ (.A1(_06496_),
    .A2(_06499_),
    .B1(net1777),
    .Y(_01700_));
 sky130_fd_sc_hd__a211o_1 _22828_ (.A1(_05527_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06478_),
    .X(_06501_));
 sky130_fd_sc_hd__nand2_1 _22829_ (.A(_06472_),
    .B(net752),
    .Y(_06502_));
 sky130_fd_sc_hd__o21ai_1 _22830_ (.A1(_06496_),
    .A2(_06501_),
    .B1(net753),
    .Y(_01701_));
 sky130_fd_sc_hd__a211o_1 _22831_ (.A1(_05530_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06481_),
    .X(_06503_));
 sky130_fd_sc_hd__nand2_1 _22832_ (.A(_06472_),
    .B(net954),
    .Y(_06504_));
 sky130_fd_sc_hd__o21ai_1 _22833_ (.A1(_06496_),
    .A2(_06503_),
    .B1(net955),
    .Y(_01702_));
 sky130_fd_sc_hd__a211o_1 _22834_ (.A1(_05533_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06484_),
    .X(_06505_));
 sky130_fd_sc_hd__nand2_1 _22835_ (.A(_06472_),
    .B(net606),
    .Y(_06506_));
 sky130_fd_sc_hd__o21ai_1 _22836_ (.A1(_06496_),
    .A2(_06505_),
    .B1(net607),
    .Y(_01703_));
 sky130_fd_sc_hd__a211o_1 _22837_ (.A1(_05536_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06487_),
    .X(_06507_));
 sky130_fd_sc_hd__nand2_1 _22838_ (.A(_06472_),
    .B(net658),
    .Y(_06508_));
 sky130_fd_sc_hd__o21ai_1 _22839_ (.A1(_06496_),
    .A2(_06507_),
    .B1(net659),
    .Y(_01704_));
 sky130_fd_sc_hd__a211o_1 _22840_ (.A1(_05539_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06490_),
    .X(_06509_));
 sky130_fd_sc_hd__nand2_1 _22841_ (.A(_06472_),
    .B(net1877),
    .Y(_06510_));
 sky130_fd_sc_hd__o21ai_1 _22842_ (.A1(_06496_),
    .A2(_06509_),
    .B1(net1878),
    .Y(_01705_));
 sky130_fd_sc_hd__a211o_1 _22843_ (.A1(_05542_),
    .A2(_06468_),
    .B1(_06477_),
    .C1(_06493_),
    .X(_06511_));
 sky130_fd_sc_hd__nand2_1 _22844_ (.A(_06472_),
    .B(net1452),
    .Y(_06512_));
 sky130_fd_sc_hd__o21ai_1 _22845_ (.A1(_06496_),
    .A2(_06511_),
    .B1(net1453),
    .Y(_01706_));
 sky130_fd_sc_hd__a211o_1 _22846_ (.A1(_05545_),
    .A2(_06469_),
    .B1(_06477_),
    .C1(_06470_),
    .X(_06513_));
 sky130_fd_sc_hd__nand2_1 _22847_ (.A(_06467_),
    .B(net1714),
    .Y(_06514_));
 sky130_fd_sc_hd__o21ai_1 _22848_ (.A1(_06496_),
    .A2(_06513_),
    .B1(net1715),
    .Y(_01707_));
 sky130_fd_sc_hd__a211o_1 _22849_ (.A1(_05548_),
    .A2(_06469_),
    .B1(_06477_),
    .C1(_06474_),
    .X(_06515_));
 sky130_fd_sc_hd__nand2_1 _22850_ (.A(_06467_),
    .B(net1044),
    .Y(_06516_));
 sky130_fd_sc_hd__o21ai_1 _22851_ (.A1(_06496_),
    .A2(_06515_),
    .B1(net1045),
    .Y(_01708_));
 sky130_fd_sc_hd__clkbuf_8 _22852_ (.A(_05892_),
    .X(_06517_));
 sky130_fd_sc_hd__a211o_1 _22853_ (.A1(_05551_),
    .A2(_06469_),
    .B1(_06517_),
    .C1(_06478_),
    .X(_06518_));
 sky130_fd_sc_hd__nand2_1 _22854_ (.A(_06467_),
    .B(net1636),
    .Y(_06519_));
 sky130_fd_sc_hd__o21ai_1 _22855_ (.A1(_06496_),
    .A2(_06518_),
    .B1(net1637),
    .Y(_01709_));
 sky130_fd_sc_hd__a211o_1 _22856_ (.A1(_05555_),
    .A2(_06469_),
    .B1(_06517_),
    .C1(_06481_),
    .X(_06520_));
 sky130_fd_sc_hd__nand2_1 _22857_ (.A(_06467_),
    .B(net1052),
    .Y(_06521_));
 sky130_fd_sc_hd__o21ai_1 _22858_ (.A1(_06496_),
    .A2(_06520_),
    .B1(net1053),
    .Y(_01710_));
 sky130_fd_sc_hd__a211o_1 _22859_ (.A1(_05558_),
    .A2(_06469_),
    .B1(_06517_),
    .C1(_06484_),
    .X(_06522_));
 sky130_fd_sc_hd__nand2_1 _22860_ (.A(_06467_),
    .B(net706),
    .Y(_06523_));
 sky130_fd_sc_hd__o21ai_1 _22861_ (.A1(_06496_),
    .A2(_06522_),
    .B1(net707),
    .Y(_01711_));
 sky130_fd_sc_hd__a211o_1 _22862_ (.A1(_05561_),
    .A2(_06469_),
    .B1(_06517_),
    .C1(_06487_),
    .X(_06524_));
 sky130_fd_sc_hd__nand2_1 _22863_ (.A(_06467_),
    .B(net1608),
    .Y(_06525_));
 sky130_fd_sc_hd__o21ai_1 _22864_ (.A1(_06496_),
    .A2(_06524_),
    .B1(net1609),
    .Y(_01712_));
 sky130_fd_sc_hd__a211o_1 _22865_ (.A1(_05564_),
    .A2(_06469_),
    .B1(_06517_),
    .C1(_06490_),
    .X(_06526_));
 sky130_fd_sc_hd__nand2_1 _22866_ (.A(_06467_),
    .B(net1316),
    .Y(_06527_));
 sky130_fd_sc_hd__o21ai_1 _22867_ (.A1(_06496_),
    .A2(_06526_),
    .B1(net1317),
    .Y(_01713_));
 sky130_fd_sc_hd__a211o_1 _22868_ (.A1(_05567_),
    .A2(_06469_),
    .B1(_06517_),
    .C1(_06493_),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_1 _22869_ (.A(_06467_),
    .B(net1296),
    .Y(_06529_));
 sky130_fd_sc_hd__o21ai_1 _22870_ (.A1(_06496_),
    .A2(_06528_),
    .B1(net1297),
    .Y(_01714_));
 sky130_fd_sc_hd__buf_8 _22871_ (.A(_02809_),
    .X(_06530_));
 sky130_fd_sc_hd__inv_2 _22872_ (.A(_12308_),
    .Y(_06531_));
 sky130_fd_sc_hd__and2_2 _22873_ (.A(_06531_),
    .B(_02813_),
    .X(_06532_));
 sky130_fd_sc_hd__nand2_1 _22874_ (.A(_06532_),
    .B(_04104_),
    .Y(_06533_));
 sky130_fd_sc_hd__buf_8 _22875_ (.A(_09109_),
    .X(_06534_));
 sky130_fd_sc_hd__a21bo_1 _22876_ (.A1(_06533_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_06535_));
 sky130_fd_sc_hd__clkbuf_8 _22877_ (.A(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__mux2_1 _22878_ (.A0(_06530_),
    .A1(net2172),
    .S(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__clkbuf_1 _22879_ (.A(_06537_),
    .X(_01715_));
 sky130_fd_sc_hd__buf_8 _22880_ (.A(_02822_),
    .X(_06538_));
 sky130_fd_sc_hd__mux2_1 _22881_ (.A0(_06538_),
    .A1(net2204),
    .S(_06536_),
    .X(_06539_));
 sky130_fd_sc_hd__clkbuf_1 _22882_ (.A(_06539_),
    .X(_01716_));
 sky130_fd_sc_hd__clkbuf_16 _22883_ (.A(_02826_),
    .X(_06540_));
 sky130_fd_sc_hd__mux2_1 _22884_ (.A0(_06540_),
    .A1(net2075),
    .S(_06536_),
    .X(_06541_));
 sky130_fd_sc_hd__clkbuf_1 _22885_ (.A(_06541_),
    .X(_01717_));
 sky130_fd_sc_hd__buf_8 _22886_ (.A(_02830_),
    .X(_06542_));
 sky130_fd_sc_hd__mux2_1 _22887_ (.A0(_06542_),
    .A1(net2136),
    .S(_06536_),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_1 _22888_ (.A(_06543_),
    .X(_01718_));
 sky130_fd_sc_hd__buf_8 _22889_ (.A(_02834_),
    .X(_06544_));
 sky130_fd_sc_hd__mux2_1 _22890_ (.A0(_06544_),
    .A1(net2295),
    .S(_06536_),
    .X(_06545_));
 sky130_fd_sc_hd__clkbuf_1 _22891_ (.A(_06545_),
    .X(_01719_));
 sky130_fd_sc_hd__clkbuf_16 _22892_ (.A(_02838_),
    .X(_06546_));
 sky130_fd_sc_hd__mux2_1 _22893_ (.A0(_06546_),
    .A1(net2525),
    .S(_06536_),
    .X(_06547_));
 sky130_fd_sc_hd__clkbuf_1 _22894_ (.A(_06547_),
    .X(_01720_));
 sky130_fd_sc_hd__buf_8 _22895_ (.A(_02842_),
    .X(_06548_));
 sky130_fd_sc_hd__mux2_1 _22896_ (.A0(_06548_),
    .A1(net2053),
    .S(_06536_),
    .X(_06549_));
 sky130_fd_sc_hd__clkbuf_1 _22897_ (.A(_06549_),
    .X(_01721_));
 sky130_fd_sc_hd__buf_8 _22898_ (.A(_02846_),
    .X(_06550_));
 sky130_fd_sc_hd__mux2_1 _22899_ (.A0(_06550_),
    .A1(net2532),
    .S(_06536_),
    .X(_06551_));
 sky130_fd_sc_hd__clkbuf_1 _22900_ (.A(_06551_),
    .X(_01722_));
 sky130_fd_sc_hd__buf_4 _22901_ (.A(_06533_),
    .X(_06552_));
 sky130_fd_sc_hd__buf_4 _22902_ (.A(_06533_),
    .X(_06553_));
 sky130_fd_sc_hd__nand2_1 _22903_ (.A(_06553_),
    .B(_05010_),
    .Y(_06554_));
 sky130_fd_sc_hd__o211a_1 _22904_ (.A1(_05095_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__mux2_1 _22905_ (.A0(_06555_),
    .A1(net2187),
    .S(_06536_),
    .X(_06556_));
 sky130_fd_sc_hd__clkbuf_1 _22906_ (.A(_06556_),
    .X(_01723_));
 sky130_fd_sc_hd__nand2_1 _22907_ (.A(_06553_),
    .B(_05014_),
    .Y(_06557_));
 sky130_fd_sc_hd__o211a_1 _22908_ (.A1(_05101_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__mux2_1 _22909_ (.A0(_06558_),
    .A1(net2381),
    .S(_06536_),
    .X(_06559_));
 sky130_fd_sc_hd__clkbuf_1 _22910_ (.A(_06559_),
    .X(_01724_));
 sky130_fd_sc_hd__nand2_1 _22911_ (.A(_06553_),
    .B(_05018_),
    .Y(_06560_));
 sky130_fd_sc_hd__o211a_1 _22912_ (.A1(_05105_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__mux2_1 _22913_ (.A0(_06561_),
    .A1(net2166),
    .S(_06536_),
    .X(_06562_));
 sky130_fd_sc_hd__clkbuf_1 _22914_ (.A(_06562_),
    .X(_01725_));
 sky130_fd_sc_hd__nand2_1 _22915_ (.A(_06553_),
    .B(_05022_),
    .Y(_06563_));
 sky130_fd_sc_hd__o211a_1 _22916_ (.A1(_05109_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__mux2_1 _22917_ (.A0(_06564_),
    .A1(net2147),
    .S(_06536_),
    .X(_06565_));
 sky130_fd_sc_hd__clkbuf_1 _22918_ (.A(_06565_),
    .X(_01726_));
 sky130_fd_sc_hd__nand2_1 _22919_ (.A(_06553_),
    .B(_05026_),
    .Y(_06566_));
 sky130_fd_sc_hd__o211a_1 _22920_ (.A1(_05113_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__mux2_1 _22921_ (.A0(_06567_),
    .A1(net2254),
    .S(_06536_),
    .X(_06568_));
 sky130_fd_sc_hd__clkbuf_1 _22922_ (.A(_06568_),
    .X(_01727_));
 sky130_fd_sc_hd__nand2_1 _22923_ (.A(_06553_),
    .B(_05030_),
    .Y(_06569_));
 sky130_fd_sc_hd__o211a_1 _22924_ (.A1(_05117_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__mux2_1 _22925_ (.A0(_06570_),
    .A1(net2049),
    .S(_06536_),
    .X(_06571_));
 sky130_fd_sc_hd__clkbuf_1 _22926_ (.A(_06571_),
    .X(_01728_));
 sky130_fd_sc_hd__nand2_1 _22927_ (.A(_06553_),
    .B(_05034_),
    .Y(_06572_));
 sky130_fd_sc_hd__o211a_1 _22928_ (.A1(_05121_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__mux2_1 _22929_ (.A0(_06573_),
    .A1(net2117),
    .S(_06536_),
    .X(_06574_));
 sky130_fd_sc_hd__clkbuf_1 _22930_ (.A(_06574_),
    .X(_01729_));
 sky130_fd_sc_hd__nand2_1 _22931_ (.A(_06553_),
    .B(_05038_),
    .Y(_06575_));
 sky130_fd_sc_hd__o211a_1 _22932_ (.A1(_05125_),
    .A2(_06552_),
    .B1(_06439_),
    .C1(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__mux2_1 _22933_ (.A0(_06576_),
    .A1(net2305),
    .S(_06536_),
    .X(_06577_));
 sky130_fd_sc_hd__clkbuf_1 _22934_ (.A(_06577_),
    .X(_01730_));
 sky130_fd_sc_hd__buf_4 _22935_ (.A(_05183_),
    .X(_06578_));
 sky130_fd_sc_hd__o211a_1 _22936_ (.A1(_05129_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06554_),
    .X(_06579_));
 sky130_fd_sc_hd__clkbuf_8 _22937_ (.A(_06535_),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _22938_ (.A0(_06579_),
    .A1(net2402),
    .S(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__clkbuf_1 _22939_ (.A(_06581_),
    .X(_01731_));
 sky130_fd_sc_hd__o211a_1 _22940_ (.A1(_05134_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06557_),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_1 _22941_ (.A0(_06582_),
    .A1(net3575),
    .S(_06580_),
    .X(_06583_));
 sky130_fd_sc_hd__clkbuf_1 _22942_ (.A(_06583_),
    .X(_01732_));
 sky130_fd_sc_hd__o211a_1 _22943_ (.A1(_05137_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06560_),
    .X(_06584_));
 sky130_fd_sc_hd__mux2_1 _22944_ (.A0(_06584_),
    .A1(net2683),
    .S(_06580_),
    .X(_06585_));
 sky130_fd_sc_hd__clkbuf_1 _22945_ (.A(_06585_),
    .X(_01733_));
 sky130_fd_sc_hd__o211a_1 _22946_ (.A1(_05140_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06563_),
    .X(_06586_));
 sky130_fd_sc_hd__mux2_1 _22947_ (.A0(_06586_),
    .A1(net2810),
    .S(_06580_),
    .X(_06587_));
 sky130_fd_sc_hd__clkbuf_1 _22948_ (.A(_06587_),
    .X(_01734_));
 sky130_fd_sc_hd__o211a_1 _22949_ (.A1(_05143_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06566_),
    .X(_06588_));
 sky130_fd_sc_hd__mux2_1 _22950_ (.A0(_06588_),
    .A1(net2669),
    .S(_06580_),
    .X(_06589_));
 sky130_fd_sc_hd__clkbuf_1 _22951_ (.A(_06589_),
    .X(_01735_));
 sky130_fd_sc_hd__o211a_1 _22952_ (.A1(_05146_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06569_),
    .X(_06590_));
 sky130_fd_sc_hd__mux2_1 _22953_ (.A0(_06590_),
    .A1(net2325),
    .S(_06580_),
    .X(_06591_));
 sky130_fd_sc_hd__clkbuf_1 _22954_ (.A(_06591_),
    .X(_01736_));
 sky130_fd_sc_hd__o211a_1 _22955_ (.A1(_05149_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06572_),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_1 _22956_ (.A0(_06592_),
    .A1(net2922),
    .S(_06580_),
    .X(_06593_));
 sky130_fd_sc_hd__clkbuf_1 _22957_ (.A(_06593_),
    .X(_01737_));
 sky130_fd_sc_hd__o211a_1 _22958_ (.A1(_05152_),
    .A2(_06552_),
    .B1(_06578_),
    .C1(_06575_),
    .X(_06594_));
 sky130_fd_sc_hd__mux2_1 _22959_ (.A0(_06594_),
    .A1(net2229),
    .S(_06580_),
    .X(_06595_));
 sky130_fd_sc_hd__clkbuf_1 _22960_ (.A(_06595_),
    .X(_01738_));
 sky130_fd_sc_hd__o211a_1 _22961_ (.A1(_05059_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06554_),
    .X(_06596_));
 sky130_fd_sc_hd__mux2_1 _22962_ (.A0(_06596_),
    .A1(net3000),
    .S(_06580_),
    .X(_06597_));
 sky130_fd_sc_hd__clkbuf_1 _22963_ (.A(_06597_),
    .X(_01739_));
 sky130_fd_sc_hd__o211a_1 _22964_ (.A1(_05063_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06557_),
    .X(_06598_));
 sky130_fd_sc_hd__mux2_1 _22965_ (.A0(_06598_),
    .A1(net3482),
    .S(_06580_),
    .X(_06599_));
 sky130_fd_sc_hd__clkbuf_1 _22966_ (.A(_06599_),
    .X(_01740_));
 sky130_fd_sc_hd__o211a_1 _22967_ (.A1(_05066_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06560_),
    .X(_06600_));
 sky130_fd_sc_hd__mux2_1 _22968_ (.A0(_06600_),
    .A1(net2615),
    .S(_06580_),
    .X(_06601_));
 sky130_fd_sc_hd__clkbuf_1 _22969_ (.A(_06601_),
    .X(_01741_));
 sky130_fd_sc_hd__o211a_1 _22970_ (.A1(_05069_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06563_),
    .X(_06602_));
 sky130_fd_sc_hd__mux2_1 _22971_ (.A0(_06602_),
    .A1(net3252),
    .S(_06580_),
    .X(_06603_));
 sky130_fd_sc_hd__clkbuf_1 _22972_ (.A(_06603_),
    .X(_01742_));
 sky130_fd_sc_hd__o211a_1 _22973_ (.A1(_05072_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06566_),
    .X(_06604_));
 sky130_fd_sc_hd__mux2_1 _22974_ (.A0(_06604_),
    .A1(net3238),
    .S(_06580_),
    .X(_06605_));
 sky130_fd_sc_hd__clkbuf_1 _22975_ (.A(_06605_),
    .X(_01743_));
 sky130_fd_sc_hd__o211a_1 _22976_ (.A1(_05075_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06569_),
    .X(_06606_));
 sky130_fd_sc_hd__mux2_1 _22977_ (.A0(_06606_),
    .A1(net2907),
    .S(_06580_),
    .X(_06607_));
 sky130_fd_sc_hd__clkbuf_1 _22978_ (.A(_06607_),
    .X(_01744_));
 sky130_fd_sc_hd__o211a_1 _22979_ (.A1(_05078_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06572_),
    .X(_06608_));
 sky130_fd_sc_hd__mux2_1 _22980_ (.A0(_06608_),
    .A1(net3102),
    .S(_06580_),
    .X(_06609_));
 sky130_fd_sc_hd__clkbuf_1 _22981_ (.A(_06609_),
    .X(_01745_));
 sky130_fd_sc_hd__o211a_1 _22982_ (.A1(_05081_),
    .A2(_06553_),
    .B1(_06578_),
    .C1(_06575_),
    .X(_06610_));
 sky130_fd_sc_hd__mux2_1 _22983_ (.A0(_06610_),
    .A1(net3035),
    .S(_06580_),
    .X(_06611_));
 sky130_fd_sc_hd__clkbuf_1 _22984_ (.A(_06611_),
    .X(_01746_));
 sky130_fd_sc_hd__nand2_1 _22985_ (.A(_06532_),
    .B(_04183_),
    .Y(_06612_));
 sky130_fd_sc_hd__a21bo_1 _22986_ (.A1(_06612_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_06613_));
 sky130_fd_sc_hd__clkbuf_8 _22987_ (.A(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__mux2_1 _22988_ (.A0(_06530_),
    .A1(net2782),
    .S(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__clkbuf_1 _22989_ (.A(_06615_),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _22990_ (.A0(_06538_),
    .A1(net3140),
    .S(_06614_),
    .X(_06616_));
 sky130_fd_sc_hd__clkbuf_1 _22991_ (.A(_06616_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _22992_ (.A0(_06540_),
    .A1(net2334),
    .S(_06614_),
    .X(_06617_));
 sky130_fd_sc_hd__clkbuf_1 _22993_ (.A(_06617_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _22994_ (.A0(_06542_),
    .A1(net2748),
    .S(_06614_),
    .X(_06618_));
 sky130_fd_sc_hd__clkbuf_1 _22995_ (.A(_06618_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _22996_ (.A0(_06544_),
    .A1(net2682),
    .S(_06614_),
    .X(_06619_));
 sky130_fd_sc_hd__clkbuf_1 _22997_ (.A(_06619_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _22998_ (.A0(_06546_),
    .A1(net3516),
    .S(_06614_),
    .X(_06620_));
 sky130_fd_sc_hd__clkbuf_1 _22999_ (.A(_06620_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _23000_ (.A0(_06548_),
    .A1(net2712),
    .S(_06614_),
    .X(_06621_));
 sky130_fd_sc_hd__clkbuf_1 _23001_ (.A(_06621_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _23002_ (.A0(_06550_),
    .A1(net2470),
    .S(_06614_),
    .X(_06622_));
 sky130_fd_sc_hd__clkbuf_1 _23003_ (.A(_06622_),
    .X(_01754_));
 sky130_fd_sc_hd__buf_4 _23004_ (.A(_06612_),
    .X(_06623_));
 sky130_fd_sc_hd__buf_4 _23005_ (.A(_05183_),
    .X(_06624_));
 sky130_fd_sc_hd__buf_4 _23006_ (.A(_06612_),
    .X(_06625_));
 sky130_fd_sc_hd__nand2_1 _23007_ (.A(_06625_),
    .B(_05010_),
    .Y(_06626_));
 sky130_fd_sc_hd__o211a_1 _23008_ (.A1(_05095_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__mux2_1 _23009_ (.A0(_06627_),
    .A1(net2419),
    .S(_06614_),
    .X(_06628_));
 sky130_fd_sc_hd__clkbuf_1 _23010_ (.A(_06628_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _23011_ (.A(_06625_),
    .B(_05014_),
    .Y(_06629_));
 sky130_fd_sc_hd__o211a_1 _23012_ (.A1(_05101_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__mux2_1 _23013_ (.A0(_06630_),
    .A1(net3236),
    .S(_06614_),
    .X(_06631_));
 sky130_fd_sc_hd__clkbuf_1 _23014_ (.A(_06631_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_1 _23015_ (.A(_06625_),
    .B(_05018_),
    .Y(_06632_));
 sky130_fd_sc_hd__o211a_1 _23016_ (.A1(_05105_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__mux2_1 _23017_ (.A0(_06633_),
    .A1(net2875),
    .S(_06614_),
    .X(_06634_));
 sky130_fd_sc_hd__clkbuf_1 _23018_ (.A(_06634_),
    .X(_01757_));
 sky130_fd_sc_hd__nand2_1 _23019_ (.A(_06625_),
    .B(_05022_),
    .Y(_06635_));
 sky130_fd_sc_hd__o211a_1 _23020_ (.A1(_05109_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__mux2_1 _23021_ (.A0(_06636_),
    .A1(net2242),
    .S(_06614_),
    .X(_06637_));
 sky130_fd_sc_hd__clkbuf_1 _23022_ (.A(_06637_),
    .X(_01758_));
 sky130_fd_sc_hd__nand2_1 _23023_ (.A(_06625_),
    .B(_05026_),
    .Y(_06638_));
 sky130_fd_sc_hd__o211a_1 _23024_ (.A1(_05113_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__mux2_1 _23025_ (.A0(_06639_),
    .A1(net3504),
    .S(_06614_),
    .X(_06640_));
 sky130_fd_sc_hd__clkbuf_1 _23026_ (.A(_06640_),
    .X(_01759_));
 sky130_fd_sc_hd__nand2_1 _23027_ (.A(_06625_),
    .B(_05030_),
    .Y(_06641_));
 sky130_fd_sc_hd__o211a_1 _23028_ (.A1(_05117_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__mux2_1 _23029_ (.A0(_06642_),
    .A1(net3369),
    .S(_06614_),
    .X(_06643_));
 sky130_fd_sc_hd__clkbuf_1 _23030_ (.A(_06643_),
    .X(_01760_));
 sky130_fd_sc_hd__nand2_1 _23031_ (.A(_06625_),
    .B(_05034_),
    .Y(_06644_));
 sky130_fd_sc_hd__o211a_1 _23032_ (.A1(_05121_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__mux2_1 _23033_ (.A0(_06645_),
    .A1(net3386),
    .S(_06614_),
    .X(_06646_));
 sky130_fd_sc_hd__clkbuf_1 _23034_ (.A(_06646_),
    .X(_01761_));
 sky130_fd_sc_hd__nand2_1 _23035_ (.A(_06625_),
    .B(_05038_),
    .Y(_06647_));
 sky130_fd_sc_hd__o211a_1 _23036_ (.A1(_05125_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__mux2_1 _23037_ (.A0(_06648_),
    .A1(net2423),
    .S(_06614_),
    .X(_06649_));
 sky130_fd_sc_hd__clkbuf_1 _23038_ (.A(_06649_),
    .X(_01762_));
 sky130_fd_sc_hd__o211a_1 _23039_ (.A1(_05129_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06626_),
    .X(_06650_));
 sky130_fd_sc_hd__clkbuf_8 _23040_ (.A(_06613_),
    .X(_06651_));
 sky130_fd_sc_hd__mux2_1 _23041_ (.A0(_06650_),
    .A1(net3336),
    .S(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__clkbuf_1 _23042_ (.A(_06652_),
    .X(_01763_));
 sky130_fd_sc_hd__o211a_1 _23043_ (.A1(_05134_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06629_),
    .X(_06653_));
 sky130_fd_sc_hd__mux2_1 _23044_ (.A0(_06653_),
    .A1(net3287),
    .S(_06651_),
    .X(_06654_));
 sky130_fd_sc_hd__clkbuf_1 _23045_ (.A(_06654_),
    .X(_01764_));
 sky130_fd_sc_hd__o211a_1 _23046_ (.A1(_05137_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06632_),
    .X(_06655_));
 sky130_fd_sc_hd__mux2_1 _23047_ (.A0(_06655_),
    .A1(net3564),
    .S(_06651_),
    .X(_06656_));
 sky130_fd_sc_hd__clkbuf_1 _23048_ (.A(_06656_),
    .X(_01765_));
 sky130_fd_sc_hd__o211a_1 _23049_ (.A1(_05140_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06635_),
    .X(_06657_));
 sky130_fd_sc_hd__mux2_1 _23050_ (.A0(_06657_),
    .A1(net2729),
    .S(_06651_),
    .X(_06658_));
 sky130_fd_sc_hd__clkbuf_1 _23051_ (.A(_06658_),
    .X(_01766_));
 sky130_fd_sc_hd__o211a_1 _23052_ (.A1(_05143_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06638_),
    .X(_06659_));
 sky130_fd_sc_hd__mux2_1 _23053_ (.A0(_06659_),
    .A1(net3589),
    .S(_06651_),
    .X(_06660_));
 sky130_fd_sc_hd__clkbuf_1 _23054_ (.A(_06660_),
    .X(_01767_));
 sky130_fd_sc_hd__o211a_1 _23055_ (.A1(_05146_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06641_),
    .X(_06661_));
 sky130_fd_sc_hd__mux2_1 _23056_ (.A0(_06661_),
    .A1(net3215),
    .S(_06651_),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_1 _23057_ (.A(_06662_),
    .X(_01768_));
 sky130_fd_sc_hd__o211a_1 _23058_ (.A1(_05149_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06644_),
    .X(_06663_));
 sky130_fd_sc_hd__mux2_1 _23059_ (.A0(_06663_),
    .A1(net3511),
    .S(_06651_),
    .X(_06664_));
 sky130_fd_sc_hd__clkbuf_1 _23060_ (.A(_06664_),
    .X(_01769_));
 sky130_fd_sc_hd__o211a_1 _23061_ (.A1(_05152_),
    .A2(_06623_),
    .B1(_06624_),
    .C1(_06647_),
    .X(_06665_));
 sky130_fd_sc_hd__mux2_1 _23062_ (.A0(_06665_),
    .A1(net3218),
    .S(_06651_),
    .X(_06666_));
 sky130_fd_sc_hd__clkbuf_1 _23063_ (.A(_06666_),
    .X(_01770_));
 sky130_fd_sc_hd__buf_4 _23064_ (.A(_05183_),
    .X(_06667_));
 sky130_fd_sc_hd__o211a_1 _23065_ (.A1(_05059_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06626_),
    .X(_06668_));
 sky130_fd_sc_hd__mux2_1 _23066_ (.A0(_06668_),
    .A1(net2426),
    .S(_06651_),
    .X(_06669_));
 sky130_fd_sc_hd__clkbuf_1 _23067_ (.A(_06669_),
    .X(_01771_));
 sky130_fd_sc_hd__o211a_1 _23068_ (.A1(_05063_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06629_),
    .X(_06670_));
 sky130_fd_sc_hd__mux2_1 _23069_ (.A0(_06670_),
    .A1(net3599),
    .S(_06651_),
    .X(_06671_));
 sky130_fd_sc_hd__clkbuf_1 _23070_ (.A(_06671_),
    .X(_01772_));
 sky130_fd_sc_hd__o211a_1 _23071_ (.A1(_05066_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06632_),
    .X(_06672_));
 sky130_fd_sc_hd__mux2_1 _23072_ (.A0(_06672_),
    .A1(net2741),
    .S(_06651_),
    .X(_06673_));
 sky130_fd_sc_hd__clkbuf_1 _23073_ (.A(_06673_),
    .X(_01773_));
 sky130_fd_sc_hd__o211a_1 _23074_ (.A1(_05069_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06635_),
    .X(_06674_));
 sky130_fd_sc_hd__mux2_1 _23075_ (.A0(_06674_),
    .A1(net2407),
    .S(_06651_),
    .X(_06675_));
 sky130_fd_sc_hd__clkbuf_1 _23076_ (.A(_06675_),
    .X(_01774_));
 sky130_fd_sc_hd__o211a_1 _23077_ (.A1(_05072_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06638_),
    .X(_06676_));
 sky130_fd_sc_hd__mux2_1 _23078_ (.A0(_06676_),
    .A1(net3552),
    .S(_06651_),
    .X(_06677_));
 sky130_fd_sc_hd__clkbuf_1 _23079_ (.A(_06677_),
    .X(_01775_));
 sky130_fd_sc_hd__o211a_1 _23080_ (.A1(_05075_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06641_),
    .X(_06678_));
 sky130_fd_sc_hd__mux2_1 _23081_ (.A0(_06678_),
    .A1(net3560),
    .S(_06651_),
    .X(_06679_));
 sky130_fd_sc_hd__clkbuf_1 _23082_ (.A(_06679_),
    .X(_01776_));
 sky130_fd_sc_hd__o211a_1 _23083_ (.A1(_05078_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06644_),
    .X(_06680_));
 sky130_fd_sc_hd__mux2_1 _23084_ (.A0(_06680_),
    .A1(net3056),
    .S(_06651_),
    .X(_06681_));
 sky130_fd_sc_hd__clkbuf_1 _23085_ (.A(_06681_),
    .X(_01777_));
 sky130_fd_sc_hd__o211a_1 _23086_ (.A1(_05081_),
    .A2(_06625_),
    .B1(_06667_),
    .C1(_06647_),
    .X(_06682_));
 sky130_fd_sc_hd__mux2_1 _23087_ (.A0(_06682_),
    .A1(net3023),
    .S(_06651_),
    .X(_06683_));
 sky130_fd_sc_hd__clkbuf_1 _23088_ (.A(_06683_),
    .X(_01778_));
 sky130_fd_sc_hd__nand2_1 _23089_ (.A(_06532_),
    .B(_04257_),
    .Y(_06684_));
 sky130_fd_sc_hd__a21bo_1 _23090_ (.A1(_06684_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_06685_));
 sky130_fd_sc_hd__clkbuf_8 _23091_ (.A(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__mux2_1 _23092_ (.A0(_06530_),
    .A1(net3445),
    .S(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__clkbuf_1 _23093_ (.A(_06687_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _23094_ (.A0(_06538_),
    .A1(net2767),
    .S(_06686_),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_1 _23095_ (.A(_06688_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _23096_ (.A0(_06540_),
    .A1(net3789),
    .S(_06686_),
    .X(_06689_));
 sky130_fd_sc_hd__clkbuf_1 _23097_ (.A(_06689_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _23098_ (.A0(_06542_),
    .A1(net2163),
    .S(_06686_),
    .X(_06690_));
 sky130_fd_sc_hd__clkbuf_1 _23099_ (.A(_06690_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _23100_ (.A0(_06544_),
    .A1(net2391),
    .S(_06686_),
    .X(_06691_));
 sky130_fd_sc_hd__clkbuf_1 _23101_ (.A(_06691_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _23102_ (.A0(_06546_),
    .A1(net2642),
    .S(_06686_),
    .X(_06692_));
 sky130_fd_sc_hd__clkbuf_1 _23103_ (.A(_06692_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _23104_ (.A0(_06548_),
    .A1(net2932),
    .S(_06686_),
    .X(_06693_));
 sky130_fd_sc_hd__clkbuf_1 _23105_ (.A(_06693_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _23106_ (.A0(_06550_),
    .A1(net2506),
    .S(_06686_),
    .X(_06694_));
 sky130_fd_sc_hd__clkbuf_1 _23107_ (.A(_06694_),
    .X(_01786_));
 sky130_fd_sc_hd__buf_4 _23108_ (.A(_06684_),
    .X(_06695_));
 sky130_fd_sc_hd__buf_4 _23109_ (.A(_06684_),
    .X(_06696_));
 sky130_fd_sc_hd__nand2_1 _23110_ (.A(_06696_),
    .B(_05010_),
    .Y(_06697_));
 sky130_fd_sc_hd__o211a_1 _23111_ (.A1(_05095_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__mux2_1 _23112_ (.A0(_06698_),
    .A1(net3078),
    .S(_06686_),
    .X(_06699_));
 sky130_fd_sc_hd__clkbuf_1 _23113_ (.A(_06699_),
    .X(_01787_));
 sky130_fd_sc_hd__nand2_1 _23114_ (.A(_06696_),
    .B(_05014_),
    .Y(_06700_));
 sky130_fd_sc_hd__o211a_1 _23115_ (.A1(_05101_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__mux2_1 _23116_ (.A0(_06701_),
    .A1(net2855),
    .S(_06686_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_1 _23117_ (.A(_06702_),
    .X(_01788_));
 sky130_fd_sc_hd__nand2_1 _23118_ (.A(_06696_),
    .B(_05018_),
    .Y(_06703_));
 sky130_fd_sc_hd__o211a_1 _23119_ (.A1(_05105_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__mux2_1 _23120_ (.A0(_06704_),
    .A1(net3199),
    .S(_06686_),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_1 _23121_ (.A(_06705_),
    .X(_01789_));
 sky130_fd_sc_hd__nand2_1 _23122_ (.A(_06696_),
    .B(_05022_),
    .Y(_06706_));
 sky130_fd_sc_hd__o211a_1 _23123_ (.A1(_05109_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__mux2_1 _23124_ (.A0(_06707_),
    .A1(net3181),
    .S(_06686_),
    .X(_06708_));
 sky130_fd_sc_hd__clkbuf_1 _23125_ (.A(_06708_),
    .X(_01790_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(_06696_),
    .B(_05026_),
    .Y(_06709_));
 sky130_fd_sc_hd__o211a_1 _23127_ (.A1(_05113_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__mux2_1 _23128_ (.A0(_06710_),
    .A1(net2699),
    .S(_06686_),
    .X(_06711_));
 sky130_fd_sc_hd__clkbuf_1 _23129_ (.A(_06711_),
    .X(_01791_));
 sky130_fd_sc_hd__nand2_1 _23130_ (.A(_06696_),
    .B(_05030_),
    .Y(_06712_));
 sky130_fd_sc_hd__o211a_1 _23131_ (.A1(_05117_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__mux2_1 _23132_ (.A0(_06713_),
    .A1(net3106),
    .S(_06686_),
    .X(_06714_));
 sky130_fd_sc_hd__clkbuf_1 _23133_ (.A(_06714_),
    .X(_01792_));
 sky130_fd_sc_hd__nand2_1 _23134_ (.A(_06696_),
    .B(_05034_),
    .Y(_06715_));
 sky130_fd_sc_hd__o211a_1 _23135_ (.A1(_05121_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__mux2_1 _23136_ (.A0(_06716_),
    .A1(net3256),
    .S(_06686_),
    .X(_06717_));
 sky130_fd_sc_hd__clkbuf_1 _23137_ (.A(_06717_),
    .X(_01793_));
 sky130_fd_sc_hd__nand2_1 _23138_ (.A(_06696_),
    .B(_05038_),
    .Y(_06718_));
 sky130_fd_sc_hd__o211a_1 _23139_ (.A1(_05125_),
    .A2(_06695_),
    .B1(_06667_),
    .C1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__mux2_1 _23140_ (.A0(_06719_),
    .A1(net2418),
    .S(_06686_),
    .X(_06720_));
 sky130_fd_sc_hd__clkbuf_1 _23141_ (.A(_06720_),
    .X(_01794_));
 sky130_fd_sc_hd__buf_4 _23142_ (.A(_05183_),
    .X(_06721_));
 sky130_fd_sc_hd__o211a_1 _23143_ (.A1(_05129_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06697_),
    .X(_06722_));
 sky130_fd_sc_hd__clkbuf_8 _23144_ (.A(_06685_),
    .X(_06723_));
 sky130_fd_sc_hd__mux2_1 _23145_ (.A0(_06722_),
    .A1(net3721),
    .S(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__clkbuf_1 _23146_ (.A(_06724_),
    .X(_01795_));
 sky130_fd_sc_hd__o211a_1 _23147_ (.A1(_05134_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06700_),
    .X(_06725_));
 sky130_fd_sc_hd__mux2_1 _23148_ (.A0(_06725_),
    .A1(net3350),
    .S(_06723_),
    .X(_06726_));
 sky130_fd_sc_hd__clkbuf_1 _23149_ (.A(_06726_),
    .X(_01796_));
 sky130_fd_sc_hd__o211a_1 _23150_ (.A1(_05137_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06703_),
    .X(_06727_));
 sky130_fd_sc_hd__mux2_1 _23151_ (.A0(_06727_),
    .A1(net2485),
    .S(_06723_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_1 _23152_ (.A(_06728_),
    .X(_01797_));
 sky130_fd_sc_hd__o211a_1 _23153_ (.A1(_05140_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06706_),
    .X(_06729_));
 sky130_fd_sc_hd__mux2_1 _23154_ (.A0(_06729_),
    .A1(net2552),
    .S(_06723_),
    .X(_06730_));
 sky130_fd_sc_hd__clkbuf_1 _23155_ (.A(_06730_),
    .X(_01798_));
 sky130_fd_sc_hd__o211a_1 _23156_ (.A1(_05143_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06709_),
    .X(_06731_));
 sky130_fd_sc_hd__mux2_1 _23157_ (.A0(_06731_),
    .A1(net3551),
    .S(_06723_),
    .X(_06732_));
 sky130_fd_sc_hd__clkbuf_1 _23158_ (.A(_06732_),
    .X(_01799_));
 sky130_fd_sc_hd__o211a_1 _23159_ (.A1(_05146_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06712_),
    .X(_06733_));
 sky130_fd_sc_hd__mux2_1 _23160_ (.A0(_06733_),
    .A1(net3651),
    .S(_06723_),
    .X(_06734_));
 sky130_fd_sc_hd__clkbuf_1 _23161_ (.A(_06734_),
    .X(_01800_));
 sky130_fd_sc_hd__o211a_1 _23162_ (.A1(_05149_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06715_),
    .X(_06735_));
 sky130_fd_sc_hd__mux2_1 _23163_ (.A0(_06735_),
    .A1(net3539),
    .S(_06723_),
    .X(_06736_));
 sky130_fd_sc_hd__clkbuf_1 _23164_ (.A(_06736_),
    .X(_01801_));
 sky130_fd_sc_hd__o211a_1 _23165_ (.A1(_05152_),
    .A2(_06695_),
    .B1(_06721_),
    .C1(_06718_),
    .X(_06737_));
 sky130_fd_sc_hd__mux2_1 _23166_ (.A0(_06737_),
    .A1(net3164),
    .S(_06723_),
    .X(_06738_));
 sky130_fd_sc_hd__clkbuf_1 _23167_ (.A(_06738_),
    .X(_01802_));
 sky130_fd_sc_hd__o211a_1 _23168_ (.A1(_05059_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06697_),
    .X(_06739_));
 sky130_fd_sc_hd__mux2_1 _23169_ (.A0(_06739_),
    .A1(net3840),
    .S(_06723_),
    .X(_06740_));
 sky130_fd_sc_hd__clkbuf_1 _23170_ (.A(_06740_),
    .X(_01803_));
 sky130_fd_sc_hd__o211a_1 _23171_ (.A1(_05063_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06700_),
    .X(_06741_));
 sky130_fd_sc_hd__mux2_1 _23172_ (.A0(_06741_),
    .A1(net3826),
    .S(_06723_),
    .X(_06742_));
 sky130_fd_sc_hd__clkbuf_1 _23173_ (.A(_06742_),
    .X(_01804_));
 sky130_fd_sc_hd__o211a_1 _23174_ (.A1(_05066_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06703_),
    .X(_06743_));
 sky130_fd_sc_hd__mux2_1 _23175_ (.A0(_06743_),
    .A1(net3062),
    .S(_06723_),
    .X(_06744_));
 sky130_fd_sc_hd__clkbuf_1 _23176_ (.A(_06744_),
    .X(_01805_));
 sky130_fd_sc_hd__o211a_1 _23177_ (.A1(_05069_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06706_),
    .X(_06745_));
 sky130_fd_sc_hd__mux2_1 _23178_ (.A0(_06745_),
    .A1(net3401),
    .S(_06723_),
    .X(_06746_));
 sky130_fd_sc_hd__clkbuf_1 _23179_ (.A(_06746_),
    .X(_01806_));
 sky130_fd_sc_hd__o211a_1 _23180_ (.A1(_05072_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06709_),
    .X(_06747_));
 sky130_fd_sc_hd__mux2_1 _23181_ (.A0(_06747_),
    .A1(net3611),
    .S(_06723_),
    .X(_06748_));
 sky130_fd_sc_hd__clkbuf_1 _23182_ (.A(_06748_),
    .X(_01807_));
 sky130_fd_sc_hd__o211a_1 _23183_ (.A1(_05075_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06712_),
    .X(_06749_));
 sky130_fd_sc_hd__mux2_1 _23184_ (.A0(_06749_),
    .A1(net3865),
    .S(_06723_),
    .X(_06750_));
 sky130_fd_sc_hd__clkbuf_1 _23185_ (.A(_06750_),
    .X(_01808_));
 sky130_fd_sc_hd__o211a_1 _23186_ (.A1(_05078_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06715_),
    .X(_06751_));
 sky130_fd_sc_hd__mux2_1 _23187_ (.A0(_06751_),
    .A1(net3687),
    .S(_06723_),
    .X(_06752_));
 sky130_fd_sc_hd__clkbuf_1 _23188_ (.A(_06752_),
    .X(_01809_));
 sky130_fd_sc_hd__o211a_1 _23189_ (.A1(_05081_),
    .A2(_06696_),
    .B1(_06721_),
    .C1(_06718_),
    .X(_06753_));
 sky130_fd_sc_hd__mux2_1 _23190_ (.A0(_06753_),
    .A1(net2263),
    .S(_06723_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_1 _23191_ (.A(_06754_),
    .X(_01810_));
 sky130_fd_sc_hd__buf_12 _23192_ (.A(_12289_),
    .X(_06755_));
 sky130_fd_sc_hd__nand2_1 _23193_ (.A(_06532_),
    .B(_04333_),
    .Y(_06756_));
 sky130_fd_sc_hd__inv_2 _23194_ (.A(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__o21ai_4 _23195_ (.A1(_06755_),
    .A2(_06757_),
    .B1(_06020_),
    .Y(_06758_));
 sky130_fd_sc_hd__mux2_1 _23196_ (.A0(_06530_),
    .A1(net2160),
    .S(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__clkbuf_1 _23197_ (.A(_06759_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _23198_ (.A0(_06538_),
    .A1(net3827),
    .S(_06758_),
    .X(_06760_));
 sky130_fd_sc_hd__clkbuf_1 _23199_ (.A(_06760_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _23200_ (.A0(_06540_),
    .A1(net2180),
    .S(_06758_),
    .X(_06761_));
 sky130_fd_sc_hd__clkbuf_1 _23201_ (.A(_06761_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _23202_ (.A0(_06542_),
    .A1(net3725),
    .S(_06758_),
    .X(_06762_));
 sky130_fd_sc_hd__clkbuf_1 _23203_ (.A(_06762_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _23204_ (.A0(_06544_),
    .A1(net3579),
    .S(_06758_),
    .X(_06763_));
 sky130_fd_sc_hd__clkbuf_1 _23205_ (.A(_06763_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _23206_ (.A0(_06546_),
    .A1(net3828),
    .S(_06758_),
    .X(_06764_));
 sky130_fd_sc_hd__clkbuf_1 _23207_ (.A(_06764_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _23208_ (.A0(_06548_),
    .A1(net2030),
    .S(_06758_),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_1 _23209_ (.A(_06765_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _23210_ (.A0(_06550_),
    .A1(net3592),
    .S(_06758_),
    .X(_06766_));
 sky130_fd_sc_hd__clkbuf_1 _23211_ (.A(_06766_),
    .X(_01818_));
 sky130_fd_sc_hd__buf_4 _23212_ (.A(_06758_),
    .X(_06767_));
 sky130_fd_sc_hd__buf_4 _23213_ (.A(_06757_),
    .X(_06768_));
 sky130_fd_sc_hd__buf_4 _23214_ (.A(_06757_),
    .X(_06769_));
 sky130_fd_sc_hd__nor2_1 _23215_ (.A(_05583_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__a211o_1 _23216_ (.A1(_05484_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__buf_4 _23217_ (.A(_06758_),
    .X(_06772_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(_06772_),
    .B(net1858),
    .Y(_06773_));
 sky130_fd_sc_hd__o21ai_1 _23219_ (.A1(_06767_),
    .A2(_06771_),
    .B1(net1859),
    .Y(_01819_));
 sky130_fd_sc_hd__nor2_1 _23220_ (.A(_05589_),
    .B(_06769_),
    .Y(_06774_));
 sky130_fd_sc_hd__a211o_1 _23221_ (.A1(_05491_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__nand2_1 _23222_ (.A(_06772_),
    .B(net1600),
    .Y(_06776_));
 sky130_fd_sc_hd__o21ai_1 _23223_ (.A1(_06767_),
    .A2(_06775_),
    .B1(net1601),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_1 _23224_ (.A(_05593_),
    .B(_06769_),
    .Y(_06777_));
 sky130_fd_sc_hd__a211o_1 _23225_ (.A1(_05495_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__nand2_1 _23226_ (.A(_06772_),
    .B(net1650),
    .Y(_06779_));
 sky130_fd_sc_hd__o21ai_1 _23227_ (.A1(_06767_),
    .A2(_06778_),
    .B1(net1651),
    .Y(_01821_));
 sky130_fd_sc_hd__nor2_1 _23228_ (.A(_05597_),
    .B(_06769_),
    .Y(_06780_));
 sky130_fd_sc_hd__a211o_1 _23229_ (.A1(_05500_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__nand2_1 _23230_ (.A(_06772_),
    .B(net1917),
    .Y(_06782_));
 sky130_fd_sc_hd__o21ai_1 _23231_ (.A1(_06767_),
    .A2(_06781_),
    .B1(net1918),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _23232_ (.A(_05601_),
    .B(_06769_),
    .Y(_06783_));
 sky130_fd_sc_hd__a211o_1 _23233_ (.A1(_05504_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__nand2_1 _23234_ (.A(_06772_),
    .B(net1244),
    .Y(_06785_));
 sky130_fd_sc_hd__o21ai_1 _23235_ (.A1(_06767_),
    .A2(_06784_),
    .B1(net1245),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _23236_ (.A(_05605_),
    .B(_06769_),
    .Y(_06786_));
 sky130_fd_sc_hd__a211o_1 _23237_ (.A1(_05508_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__nand2_1 _23238_ (.A(_06772_),
    .B(net1720),
    .Y(_06788_));
 sky130_fd_sc_hd__o21ai_1 _23239_ (.A1(_06767_),
    .A2(_06787_),
    .B1(net1721),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _23240_ (.A(_05609_),
    .B(_06769_),
    .Y(_06789_));
 sky130_fd_sc_hd__a211o_1 _23241_ (.A1(_05512_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__nand2_1 _23242_ (.A(_06772_),
    .B(net1956),
    .Y(_06791_));
 sky130_fd_sc_hd__o21ai_1 _23243_ (.A1(_06767_),
    .A2(_06790_),
    .B1(net1957),
    .Y(_01825_));
 sky130_fd_sc_hd__nor2_1 _23244_ (.A(_05613_),
    .B(_06769_),
    .Y(_06792_));
 sky130_fd_sc_hd__a211o_1 _23245_ (.A1(_05516_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_1 _23246_ (.A(_06772_),
    .B(net1628),
    .Y(_06794_));
 sky130_fd_sc_hd__o21ai_1 _23247_ (.A1(_06767_),
    .A2(_06793_),
    .B1(net1629),
    .Y(_01826_));
 sky130_fd_sc_hd__buf_4 _23248_ (.A(_06758_),
    .X(_06795_));
 sky130_fd_sc_hd__a211o_1 _23249_ (.A1(_05521_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06770_),
    .X(_06796_));
 sky130_fd_sc_hd__nand2_1 _23250_ (.A(_06772_),
    .B(net1604),
    .Y(_06797_));
 sky130_fd_sc_hd__o21ai_1 _23251_ (.A1(_06795_),
    .A2(_06796_),
    .B1(net1605),
    .Y(_01827_));
 sky130_fd_sc_hd__a211o_1 _23252_ (.A1(_05524_),
    .A2(_06768_),
    .B1(_06517_),
    .C1(_06774_),
    .X(_06798_));
 sky130_fd_sc_hd__nand2_1 _23253_ (.A(_06772_),
    .B(net1810),
    .Y(_06799_));
 sky130_fd_sc_hd__o21ai_1 _23254_ (.A1(_06795_),
    .A2(_06798_),
    .B1(net1811),
    .Y(_01828_));
 sky130_fd_sc_hd__buf_4 _23255_ (.A(_05892_),
    .X(_06800_));
 sky130_fd_sc_hd__a211o_1 _23256_ (.A1(_05527_),
    .A2(_06768_),
    .B1(_06800_),
    .C1(_06777_),
    .X(_06801_));
 sky130_fd_sc_hd__nand2_1 _23257_ (.A(_06772_),
    .B(net1166),
    .Y(_06802_));
 sky130_fd_sc_hd__o21ai_1 _23258_ (.A1(_06795_),
    .A2(_06801_),
    .B1(net1167),
    .Y(_01829_));
 sky130_fd_sc_hd__a211o_1 _23259_ (.A1(_05530_),
    .A2(_06768_),
    .B1(_06800_),
    .C1(_06780_),
    .X(_06803_));
 sky130_fd_sc_hd__nand2_1 _23260_ (.A(_06772_),
    .B(net1915),
    .Y(_06804_));
 sky130_fd_sc_hd__o21ai_1 _23261_ (.A1(_06795_),
    .A2(_06803_),
    .B1(net1916),
    .Y(_01830_));
 sky130_fd_sc_hd__a211o_1 _23262_ (.A1(_05533_),
    .A2(_06768_),
    .B1(_06800_),
    .C1(_06783_),
    .X(_06805_));
 sky130_fd_sc_hd__nand2_1 _23263_ (.A(_06772_),
    .B(net1274),
    .Y(_06806_));
 sky130_fd_sc_hd__o21ai_1 _23264_ (.A1(_06795_),
    .A2(_06805_),
    .B1(net1275),
    .Y(_01831_));
 sky130_fd_sc_hd__a211o_1 _23265_ (.A1(_05536_),
    .A2(_06768_),
    .B1(_06800_),
    .C1(_06786_),
    .X(_06807_));
 sky130_fd_sc_hd__nand2_1 _23266_ (.A(_06772_),
    .B(net750),
    .Y(_06808_));
 sky130_fd_sc_hd__o21ai_1 _23267_ (.A1(_06795_),
    .A2(_06807_),
    .B1(net751),
    .Y(_01832_));
 sky130_fd_sc_hd__a211o_1 _23268_ (.A1(_05539_),
    .A2(_06768_),
    .B1(_06800_),
    .C1(_06789_),
    .X(_06809_));
 sky130_fd_sc_hd__nand2_1 _23269_ (.A(_06772_),
    .B(net1396),
    .Y(_06810_));
 sky130_fd_sc_hd__o21ai_1 _23270_ (.A1(_06795_),
    .A2(_06809_),
    .B1(net1397),
    .Y(_01833_));
 sky130_fd_sc_hd__a211o_1 _23271_ (.A1(_05542_),
    .A2(_06768_),
    .B1(_06800_),
    .C1(_06792_),
    .X(_06811_));
 sky130_fd_sc_hd__nand2_1 _23272_ (.A(_06772_),
    .B(net1766),
    .Y(_06812_));
 sky130_fd_sc_hd__o21ai_1 _23273_ (.A1(_06795_),
    .A2(_06811_),
    .B1(net1767),
    .Y(_01834_));
 sky130_fd_sc_hd__a211o_1 _23274_ (.A1(_05545_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06770_),
    .X(_06813_));
 sky130_fd_sc_hd__nand2_1 _23275_ (.A(_06767_),
    .B(net1602),
    .Y(_06814_));
 sky130_fd_sc_hd__o21ai_1 _23276_ (.A1(_06795_),
    .A2(_06813_),
    .B1(net1603),
    .Y(_01835_));
 sky130_fd_sc_hd__a211o_1 _23277_ (.A1(_05548_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06774_),
    .X(_06815_));
 sky130_fd_sc_hd__nand2_1 _23278_ (.A(_06767_),
    .B(net1963),
    .Y(_06816_));
 sky130_fd_sc_hd__o21ai_1 _23279_ (.A1(_06795_),
    .A2(_06815_),
    .B1(_06816_),
    .Y(_01836_));
 sky130_fd_sc_hd__a211o_1 _23280_ (.A1(_05551_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06777_),
    .X(_06817_));
 sky130_fd_sc_hd__nand2_1 _23281_ (.A(_06767_),
    .B(net2002),
    .Y(_06818_));
 sky130_fd_sc_hd__o21ai_1 _23282_ (.A1(_06795_),
    .A2(_06817_),
    .B1(_06818_),
    .Y(_01837_));
 sky130_fd_sc_hd__a211o_1 _23283_ (.A1(_05555_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06780_),
    .X(_06819_));
 sky130_fd_sc_hd__nand2_1 _23284_ (.A(_06767_),
    .B(net1116),
    .Y(_06820_));
 sky130_fd_sc_hd__o21ai_1 _23285_ (.A1(_06795_),
    .A2(_06819_),
    .B1(net1117),
    .Y(_01838_));
 sky130_fd_sc_hd__a211o_1 _23286_ (.A1(_05558_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06783_),
    .X(_06821_));
 sky130_fd_sc_hd__nand2_1 _23287_ (.A(_06767_),
    .B(net1560),
    .Y(_06822_));
 sky130_fd_sc_hd__o21ai_1 _23288_ (.A1(_06795_),
    .A2(_06821_),
    .B1(net1561),
    .Y(_01839_));
 sky130_fd_sc_hd__a211o_1 _23289_ (.A1(_05561_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06786_),
    .X(_06823_));
 sky130_fd_sc_hd__nand2_1 _23290_ (.A(_06767_),
    .B(net786),
    .Y(_06824_));
 sky130_fd_sc_hd__o21ai_1 _23291_ (.A1(_06795_),
    .A2(_06823_),
    .B1(net787),
    .Y(_01840_));
 sky130_fd_sc_hd__a211o_1 _23292_ (.A1(_05564_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06789_),
    .X(_06825_));
 sky130_fd_sc_hd__nand2_1 _23293_ (.A(_06767_),
    .B(net936),
    .Y(_06826_));
 sky130_fd_sc_hd__o21ai_1 _23294_ (.A1(_06795_),
    .A2(_06825_),
    .B1(net937),
    .Y(_01841_));
 sky130_fd_sc_hd__a211o_1 _23295_ (.A1(_05567_),
    .A2(_06769_),
    .B1(_06800_),
    .C1(_06792_),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_1 _23296_ (.A(_06767_),
    .B(net1806),
    .Y(_06828_));
 sky130_fd_sc_hd__o21ai_1 _23297_ (.A1(_06795_),
    .A2(_06827_),
    .B1(net1807),
    .Y(_01842_));
 sky130_fd_sc_hd__and2_2 _23298_ (.A(_03207_),
    .B(_06531_),
    .X(_06829_));
 sky130_fd_sc_hd__nand2_1 _23299_ (.A(_06829_),
    .B(_04104_),
    .Y(_06830_));
 sky130_fd_sc_hd__a21bo_1 _23300_ (.A1(_06830_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_06831_));
 sky130_fd_sc_hd__clkbuf_8 _23301_ (.A(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__mux2_1 _23302_ (.A0(_06530_),
    .A1(net3666),
    .S(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__clkbuf_1 _23303_ (.A(_06833_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _23304_ (.A0(_06538_),
    .A1(net3419),
    .S(_06832_),
    .X(_06834_));
 sky130_fd_sc_hd__clkbuf_1 _23305_ (.A(_06834_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _23306_ (.A0(_06540_),
    .A1(net3095),
    .S(_06832_),
    .X(_06835_));
 sky130_fd_sc_hd__clkbuf_1 _23307_ (.A(_06835_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _23308_ (.A0(_06542_),
    .A1(net2244),
    .S(_06832_),
    .X(_06836_));
 sky130_fd_sc_hd__clkbuf_1 _23309_ (.A(_06836_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _23310_ (.A0(_06544_),
    .A1(net2328),
    .S(_06832_),
    .X(_06837_));
 sky130_fd_sc_hd__clkbuf_1 _23311_ (.A(_06837_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _23312_ (.A0(_06546_),
    .A1(net3179),
    .S(_06832_),
    .X(_06838_));
 sky130_fd_sc_hd__clkbuf_1 _23313_ (.A(_06838_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _23314_ (.A0(_06548_),
    .A1(net2197),
    .S(_06832_),
    .X(_06839_));
 sky130_fd_sc_hd__clkbuf_1 _23315_ (.A(_06839_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _23316_ (.A0(_06550_),
    .A1(net2287),
    .S(_06832_),
    .X(_06840_));
 sky130_fd_sc_hd__clkbuf_1 _23317_ (.A(_06840_),
    .X(_01850_));
 sky130_fd_sc_hd__buf_4 _23318_ (.A(_06830_),
    .X(_06841_));
 sky130_fd_sc_hd__buf_4 _23319_ (.A(_05183_),
    .X(_06842_));
 sky130_fd_sc_hd__buf_4 _23320_ (.A(_06830_),
    .X(_06843_));
 sky130_fd_sc_hd__nand2_1 _23321_ (.A(_06843_),
    .B(_05010_),
    .Y(_06844_));
 sky130_fd_sc_hd__o211a_1 _23322_ (.A1(_05095_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__mux2_1 _23323_ (.A0(_06845_),
    .A1(net3734),
    .S(_06832_),
    .X(_06846_));
 sky130_fd_sc_hd__clkbuf_1 _23324_ (.A(_06846_),
    .X(_01851_));
 sky130_fd_sc_hd__nand2_1 _23325_ (.A(_06843_),
    .B(_05014_),
    .Y(_06847_));
 sky130_fd_sc_hd__o211a_1 _23326_ (.A1(_05101_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__mux2_1 _23327_ (.A0(_06848_),
    .A1(net2820),
    .S(_06832_),
    .X(_06849_));
 sky130_fd_sc_hd__clkbuf_1 _23328_ (.A(_06849_),
    .X(_01852_));
 sky130_fd_sc_hd__nand2_1 _23329_ (.A(_06843_),
    .B(_05018_),
    .Y(_06850_));
 sky130_fd_sc_hd__o211a_1 _23330_ (.A1(_05105_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__mux2_1 _23331_ (.A0(_06851_),
    .A1(net2716),
    .S(_06832_),
    .X(_06852_));
 sky130_fd_sc_hd__clkbuf_1 _23332_ (.A(_06852_),
    .X(_01853_));
 sky130_fd_sc_hd__nand2_1 _23333_ (.A(_06843_),
    .B(_05022_),
    .Y(_06853_));
 sky130_fd_sc_hd__o211a_1 _23334_ (.A1(_05109_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__mux2_1 _23335_ (.A0(_06854_),
    .A1(net2408),
    .S(_06832_),
    .X(_06855_));
 sky130_fd_sc_hd__clkbuf_1 _23336_ (.A(_06855_),
    .X(_01854_));
 sky130_fd_sc_hd__nand2_1 _23337_ (.A(_06843_),
    .B(_05026_),
    .Y(_06856_));
 sky130_fd_sc_hd__o211a_1 _23338_ (.A1(_05113_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__mux2_1 _23339_ (.A0(_06857_),
    .A1(net3366),
    .S(_06832_),
    .X(_06858_));
 sky130_fd_sc_hd__clkbuf_1 _23340_ (.A(_06858_),
    .X(_01855_));
 sky130_fd_sc_hd__nand2_1 _23341_ (.A(_06843_),
    .B(_05030_),
    .Y(_06859_));
 sky130_fd_sc_hd__o211a_1 _23342_ (.A1(_05117_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__mux2_1 _23343_ (.A0(_06860_),
    .A1(net3493),
    .S(_06832_),
    .X(_06861_));
 sky130_fd_sc_hd__clkbuf_1 _23344_ (.A(_06861_),
    .X(_01856_));
 sky130_fd_sc_hd__nand2_1 _23345_ (.A(_06843_),
    .B(_05034_),
    .Y(_06862_));
 sky130_fd_sc_hd__o211a_1 _23346_ (.A1(_05121_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__mux2_1 _23347_ (.A0(_06863_),
    .A1(net2861),
    .S(_06832_),
    .X(_06864_));
 sky130_fd_sc_hd__clkbuf_1 _23348_ (.A(_06864_),
    .X(_01857_));
 sky130_fd_sc_hd__nand2_1 _23349_ (.A(_06843_),
    .B(_05038_),
    .Y(_06865_));
 sky130_fd_sc_hd__o211a_1 _23350_ (.A1(_05125_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06865_),
    .X(_06866_));
 sky130_fd_sc_hd__mux2_1 _23351_ (.A0(_06866_),
    .A1(net2867),
    .S(_06832_),
    .X(_06867_));
 sky130_fd_sc_hd__clkbuf_1 _23352_ (.A(_06867_),
    .X(_01858_));
 sky130_fd_sc_hd__o211a_1 _23353_ (.A1(_05129_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06844_),
    .X(_06868_));
 sky130_fd_sc_hd__clkbuf_8 _23354_ (.A(_06831_),
    .X(_06869_));
 sky130_fd_sc_hd__mux2_1 _23355_ (.A0(_06868_),
    .A1(net3724),
    .S(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__clkbuf_1 _23356_ (.A(_06870_),
    .X(_01859_));
 sky130_fd_sc_hd__o211a_1 _23357_ (.A1(_05134_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06847_),
    .X(_06871_));
 sky130_fd_sc_hd__mux2_1 _23358_ (.A0(_06871_),
    .A1(net3727),
    .S(_06869_),
    .X(_06872_));
 sky130_fd_sc_hd__clkbuf_1 _23359_ (.A(_06872_),
    .X(_01860_));
 sky130_fd_sc_hd__o211a_1 _23360_ (.A1(_05137_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06850_),
    .X(_06873_));
 sky130_fd_sc_hd__mux2_1 _23361_ (.A0(_06873_),
    .A1(net3395),
    .S(_06869_),
    .X(_06874_));
 sky130_fd_sc_hd__clkbuf_1 _23362_ (.A(_06874_),
    .X(_01861_));
 sky130_fd_sc_hd__o211a_1 _23363_ (.A1(_05140_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06853_),
    .X(_06875_));
 sky130_fd_sc_hd__mux2_1 _23364_ (.A0(_06875_),
    .A1(net3163),
    .S(_06869_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_1 _23365_ (.A(_06876_),
    .X(_01862_));
 sky130_fd_sc_hd__o211a_1 _23366_ (.A1(_05143_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06856_),
    .X(_06877_));
 sky130_fd_sc_hd__mux2_1 _23367_ (.A0(_06877_),
    .A1(net3574),
    .S(_06869_),
    .X(_06878_));
 sky130_fd_sc_hd__clkbuf_1 _23368_ (.A(_06878_),
    .X(_01863_));
 sky130_fd_sc_hd__o211a_1 _23369_ (.A1(_05146_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06859_),
    .X(_06879_));
 sky130_fd_sc_hd__mux2_1 _23370_ (.A0(_06879_),
    .A1(net2951),
    .S(_06869_),
    .X(_06880_));
 sky130_fd_sc_hd__clkbuf_1 _23371_ (.A(_06880_),
    .X(_01864_));
 sky130_fd_sc_hd__o211a_1 _23372_ (.A1(_05149_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06862_),
    .X(_06881_));
 sky130_fd_sc_hd__mux2_1 _23373_ (.A0(_06881_),
    .A1(net3282),
    .S(_06869_),
    .X(_06882_));
 sky130_fd_sc_hd__clkbuf_1 _23374_ (.A(_06882_),
    .X(_01865_));
 sky130_fd_sc_hd__o211a_1 _23375_ (.A1(_05152_),
    .A2(_06841_),
    .B1(_06842_),
    .C1(_06865_),
    .X(_06883_));
 sky130_fd_sc_hd__mux2_1 _23376_ (.A0(_06883_),
    .A1(net3143),
    .S(_06869_),
    .X(_06884_));
 sky130_fd_sc_hd__clkbuf_1 _23377_ (.A(_06884_),
    .X(_01866_));
 sky130_fd_sc_hd__buf_8 _23378_ (.A(net49),
    .X(_06885_));
 sky130_fd_sc_hd__buf_4 _23379_ (.A(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__o211a_1 _23380_ (.A1(_05059_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06844_),
    .X(_06887_));
 sky130_fd_sc_hd__mux2_1 _23381_ (.A0(_06887_),
    .A1(net2354),
    .S(_06869_),
    .X(_06888_));
 sky130_fd_sc_hd__clkbuf_1 _23382_ (.A(_06888_),
    .X(_01867_));
 sky130_fd_sc_hd__o211a_1 _23383_ (.A1(_05063_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06847_),
    .X(_06889_));
 sky130_fd_sc_hd__mux2_1 _23384_ (.A0(_06889_),
    .A1(net3276),
    .S(_06869_),
    .X(_06890_));
 sky130_fd_sc_hd__clkbuf_1 _23385_ (.A(_06890_),
    .X(_01868_));
 sky130_fd_sc_hd__o211a_1 _23386_ (.A1(_05066_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06850_),
    .X(_06891_));
 sky130_fd_sc_hd__mux2_1 _23387_ (.A0(_06891_),
    .A1(net2087),
    .S(_06869_),
    .X(_06892_));
 sky130_fd_sc_hd__clkbuf_1 _23388_ (.A(_06892_),
    .X(_01869_));
 sky130_fd_sc_hd__o211a_1 _23389_ (.A1(_05069_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06853_),
    .X(_06893_));
 sky130_fd_sc_hd__mux2_1 _23390_ (.A0(_06893_),
    .A1(net2092),
    .S(_06869_),
    .X(_06894_));
 sky130_fd_sc_hd__clkbuf_1 _23391_ (.A(_06894_),
    .X(_01870_));
 sky130_fd_sc_hd__o211a_1 _23392_ (.A1(_05072_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06856_),
    .X(_06895_));
 sky130_fd_sc_hd__mux2_1 _23393_ (.A0(_06895_),
    .A1(net3012),
    .S(_06869_),
    .X(_06896_));
 sky130_fd_sc_hd__clkbuf_1 _23394_ (.A(_06896_),
    .X(_01871_));
 sky130_fd_sc_hd__o211a_1 _23395_ (.A1(_05075_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06859_),
    .X(_06897_));
 sky130_fd_sc_hd__mux2_1 _23396_ (.A0(_06897_),
    .A1(net2102),
    .S(_06869_),
    .X(_06898_));
 sky130_fd_sc_hd__clkbuf_1 _23397_ (.A(_06898_),
    .X(_01872_));
 sky130_fd_sc_hd__o211a_1 _23398_ (.A1(_05078_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06862_),
    .X(_06899_));
 sky130_fd_sc_hd__mux2_1 _23399_ (.A0(_06899_),
    .A1(net2073),
    .S(_06869_),
    .X(_06900_));
 sky130_fd_sc_hd__clkbuf_1 _23400_ (.A(_06900_),
    .X(_01873_));
 sky130_fd_sc_hd__o211a_1 _23401_ (.A1(_05081_),
    .A2(_06843_),
    .B1(_06886_),
    .C1(_06865_),
    .X(_06901_));
 sky130_fd_sc_hd__mux2_1 _23402_ (.A0(_06901_),
    .A1(net2134),
    .S(_06869_),
    .X(_06902_));
 sky130_fd_sc_hd__clkbuf_1 _23403_ (.A(_06902_),
    .X(_01874_));
 sky130_fd_sc_hd__nand2_1 _23404_ (.A(_06829_),
    .B(_04183_),
    .Y(_06903_));
 sky130_fd_sc_hd__a21bo_1 _23405_ (.A1(_06903_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_06904_));
 sky130_fd_sc_hd__clkbuf_8 _23406_ (.A(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__mux2_1 _23407_ (.A0(_06530_),
    .A1(net2063),
    .S(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__clkbuf_1 _23408_ (.A(_06906_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _23409_ (.A0(_06538_),
    .A1(net2194),
    .S(_06905_),
    .X(_06907_));
 sky130_fd_sc_hd__clkbuf_1 _23410_ (.A(_06907_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _23411_ (.A0(_06540_),
    .A1(net2038),
    .S(_06905_),
    .X(_06908_));
 sky130_fd_sc_hd__clkbuf_1 _23412_ (.A(_06908_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _23413_ (.A0(_06542_),
    .A1(net2121),
    .S(_06905_),
    .X(_06909_));
 sky130_fd_sc_hd__clkbuf_1 _23414_ (.A(_06909_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _23415_ (.A0(_06544_),
    .A1(net2668),
    .S(_06905_),
    .X(_06910_));
 sky130_fd_sc_hd__clkbuf_1 _23416_ (.A(_06910_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _23417_ (.A0(_06546_),
    .A1(net2173),
    .S(_06905_),
    .X(_06911_));
 sky130_fd_sc_hd__clkbuf_1 _23418_ (.A(_06911_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _23419_ (.A0(_06548_),
    .A1(net2042),
    .S(_06905_),
    .X(_06912_));
 sky130_fd_sc_hd__clkbuf_1 _23420_ (.A(_06912_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _23421_ (.A0(_06550_),
    .A1(net2125),
    .S(_06905_),
    .X(_06913_));
 sky130_fd_sc_hd__clkbuf_1 _23422_ (.A(_06913_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_4 _23423_ (.A(_06903_),
    .X(_06914_));
 sky130_fd_sc_hd__buf_4 _23424_ (.A(_06903_),
    .X(_06915_));
 sky130_fd_sc_hd__nand2_1 _23425_ (.A(_06915_),
    .B(_05010_),
    .Y(_06916_));
 sky130_fd_sc_hd__o211a_1 _23426_ (.A1(_05095_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__mux2_1 _23427_ (.A0(_06917_),
    .A1(net2141),
    .S(_06905_),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_1 _23428_ (.A(_06918_),
    .X(_01883_));
 sky130_fd_sc_hd__nand2_1 _23429_ (.A(_06915_),
    .B(_05014_),
    .Y(_06919_));
 sky130_fd_sc_hd__o211a_1 _23430_ (.A1(_05101_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__mux2_1 _23431_ (.A0(_06920_),
    .A1(net3362),
    .S(_06905_),
    .X(_06921_));
 sky130_fd_sc_hd__clkbuf_1 _23432_ (.A(_06921_),
    .X(_01884_));
 sky130_fd_sc_hd__nand2_1 _23433_ (.A(_06915_),
    .B(_05018_),
    .Y(_06922_));
 sky130_fd_sc_hd__o211a_1 _23434_ (.A1(_05105_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__mux2_1 _23435_ (.A0(_06923_),
    .A1(net3585),
    .S(_06905_),
    .X(_06924_));
 sky130_fd_sc_hd__clkbuf_1 _23436_ (.A(_06924_),
    .X(_01885_));
 sky130_fd_sc_hd__nand2_1 _23437_ (.A(_06915_),
    .B(_05022_),
    .Y(_06925_));
 sky130_fd_sc_hd__o211a_1 _23438_ (.A1(_05109_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__mux2_1 _23439_ (.A0(_06926_),
    .A1(net2145),
    .S(_06905_),
    .X(_06927_));
 sky130_fd_sc_hd__clkbuf_1 _23440_ (.A(_06927_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_1 _23441_ (.A(_06915_),
    .B(_05026_),
    .Y(_06928_));
 sky130_fd_sc_hd__o211a_1 _23442_ (.A1(_05113_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__mux2_1 _23443_ (.A0(_06929_),
    .A1(net2146),
    .S(_06905_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_1 _23444_ (.A(_06930_),
    .X(_01887_));
 sky130_fd_sc_hd__nand2_1 _23445_ (.A(_06915_),
    .B(_05030_),
    .Y(_06931_));
 sky130_fd_sc_hd__o211a_1 _23446_ (.A1(_05117_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__mux2_1 _23447_ (.A0(_06932_),
    .A1(net2070),
    .S(_06905_),
    .X(_06933_));
 sky130_fd_sc_hd__clkbuf_1 _23448_ (.A(_06933_),
    .X(_01888_));
 sky130_fd_sc_hd__nand2_1 _23449_ (.A(_06915_),
    .B(_05034_),
    .Y(_06934_));
 sky130_fd_sc_hd__o211a_1 _23450_ (.A1(_05121_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__mux2_1 _23451_ (.A0(_06935_),
    .A1(net2085),
    .S(_06905_),
    .X(_06936_));
 sky130_fd_sc_hd__clkbuf_1 _23452_ (.A(_06936_),
    .X(_01889_));
 sky130_fd_sc_hd__nand2_1 _23453_ (.A(_06915_),
    .B(_05038_),
    .Y(_06937_));
 sky130_fd_sc_hd__o211a_1 _23454_ (.A1(_05125_),
    .A2(_06914_),
    .B1(_06886_),
    .C1(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__mux2_1 _23455_ (.A0(_06938_),
    .A1(net2710),
    .S(_06905_),
    .X(_06939_));
 sky130_fd_sc_hd__clkbuf_1 _23456_ (.A(_06939_),
    .X(_01890_));
 sky130_fd_sc_hd__buf_4 _23457_ (.A(_06885_),
    .X(_06940_));
 sky130_fd_sc_hd__o211a_1 _23458_ (.A1(_05129_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06916_),
    .X(_06941_));
 sky130_fd_sc_hd__clkbuf_8 _23459_ (.A(_06904_),
    .X(_06942_));
 sky130_fd_sc_hd__mux2_1 _23460_ (.A0(_06941_),
    .A1(net2378),
    .S(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__clkbuf_1 _23461_ (.A(_06943_),
    .X(_01891_));
 sky130_fd_sc_hd__o211a_1 _23462_ (.A1(_05134_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06919_),
    .X(_06944_));
 sky130_fd_sc_hd__mux2_1 _23463_ (.A0(_06944_),
    .A1(net3423),
    .S(_06942_),
    .X(_06945_));
 sky130_fd_sc_hd__clkbuf_1 _23464_ (.A(_06945_),
    .X(_01892_));
 sky130_fd_sc_hd__o211a_1 _23465_ (.A1(_05137_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06922_),
    .X(_06946_));
 sky130_fd_sc_hd__mux2_1 _23466_ (.A0(_06946_),
    .A1(net3459),
    .S(_06942_),
    .X(_06947_));
 sky130_fd_sc_hd__clkbuf_1 _23467_ (.A(_06947_),
    .X(_01893_));
 sky130_fd_sc_hd__o211a_1 _23468_ (.A1(_05140_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06925_),
    .X(_06948_));
 sky130_fd_sc_hd__mux2_1 _23469_ (.A0(_06948_),
    .A1(net2529),
    .S(_06942_),
    .X(_06949_));
 sky130_fd_sc_hd__clkbuf_1 _23470_ (.A(_06949_),
    .X(_01894_));
 sky130_fd_sc_hd__o211a_1 _23471_ (.A1(_05143_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06928_),
    .X(_06950_));
 sky130_fd_sc_hd__mux2_1 _23472_ (.A0(_06950_),
    .A1(net2065),
    .S(_06942_),
    .X(_06951_));
 sky130_fd_sc_hd__clkbuf_1 _23473_ (.A(_06951_),
    .X(_01895_));
 sky130_fd_sc_hd__o211a_1 _23474_ (.A1(_05146_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06931_),
    .X(_06952_));
 sky130_fd_sc_hd__mux2_1 _23475_ (.A0(_06952_),
    .A1(net2076),
    .S(_06942_),
    .X(_06953_));
 sky130_fd_sc_hd__clkbuf_1 _23476_ (.A(_06953_),
    .X(_01896_));
 sky130_fd_sc_hd__o211a_1 _23477_ (.A1(_05149_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06934_),
    .X(_06954_));
 sky130_fd_sc_hd__mux2_1 _23478_ (.A0(_06954_),
    .A1(net2435),
    .S(_06942_),
    .X(_06955_));
 sky130_fd_sc_hd__clkbuf_1 _23479_ (.A(_06955_),
    .X(_01897_));
 sky130_fd_sc_hd__o211a_1 _23480_ (.A1(_05152_),
    .A2(_06914_),
    .B1(_06940_),
    .C1(_06937_),
    .X(_06956_));
 sky130_fd_sc_hd__mux2_1 _23481_ (.A0(_06956_),
    .A1(net2061),
    .S(_06942_),
    .X(_06957_));
 sky130_fd_sc_hd__clkbuf_1 _23482_ (.A(_06957_),
    .X(_01898_));
 sky130_fd_sc_hd__o211a_1 _23483_ (.A1(_05059_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06916_),
    .X(_06958_));
 sky130_fd_sc_hd__mux2_1 _23484_ (.A0(_06958_),
    .A1(net3132),
    .S(_06942_),
    .X(_06959_));
 sky130_fd_sc_hd__clkbuf_1 _23485_ (.A(_06959_),
    .X(_01899_));
 sky130_fd_sc_hd__o211a_1 _23486_ (.A1(_05063_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06919_),
    .X(_06960_));
 sky130_fd_sc_hd__mux2_1 _23487_ (.A0(_06960_),
    .A1(net3739),
    .S(_06942_),
    .X(_06961_));
 sky130_fd_sc_hd__clkbuf_1 _23488_ (.A(_06961_),
    .X(_01900_));
 sky130_fd_sc_hd__o211a_1 _23489_ (.A1(_05066_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06922_),
    .X(_06962_));
 sky130_fd_sc_hd__mux2_1 _23490_ (.A0(_06962_),
    .A1(net3803),
    .S(_06942_),
    .X(_06963_));
 sky130_fd_sc_hd__clkbuf_1 _23491_ (.A(_06963_),
    .X(_01901_));
 sky130_fd_sc_hd__o211a_1 _23492_ (.A1(_05069_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06925_),
    .X(_06964_));
 sky130_fd_sc_hd__mux2_1 _23493_ (.A0(_06964_),
    .A1(net3629),
    .S(_06942_),
    .X(_06965_));
 sky130_fd_sc_hd__clkbuf_1 _23494_ (.A(_06965_),
    .X(_01902_));
 sky130_fd_sc_hd__o211a_1 _23495_ (.A1(_05072_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06928_),
    .X(_06966_));
 sky130_fd_sc_hd__mux2_1 _23496_ (.A0(_06966_),
    .A1(net3759),
    .S(_06942_),
    .X(_06967_));
 sky130_fd_sc_hd__clkbuf_1 _23497_ (.A(_06967_),
    .X(_01903_));
 sky130_fd_sc_hd__o211a_1 _23498_ (.A1(_05075_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06931_),
    .X(_06968_));
 sky130_fd_sc_hd__mux2_1 _23499_ (.A0(_06968_),
    .A1(net3744),
    .S(_06942_),
    .X(_06969_));
 sky130_fd_sc_hd__clkbuf_1 _23500_ (.A(_06969_),
    .X(_01904_));
 sky130_fd_sc_hd__o211a_1 _23501_ (.A1(_05078_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06934_),
    .X(_06970_));
 sky130_fd_sc_hd__mux2_1 _23502_ (.A0(_06970_),
    .A1(net3598),
    .S(_06942_),
    .X(_06971_));
 sky130_fd_sc_hd__clkbuf_1 _23503_ (.A(_06971_),
    .X(_01905_));
 sky130_fd_sc_hd__o211a_1 _23504_ (.A1(_05081_),
    .A2(_06915_),
    .B1(_06940_),
    .C1(_06937_),
    .X(_06972_));
 sky130_fd_sc_hd__mux2_1 _23505_ (.A0(_06972_),
    .A1(net3021),
    .S(_06942_),
    .X(_06973_));
 sky130_fd_sc_hd__clkbuf_1 _23506_ (.A(_06973_),
    .X(_01906_));
 sky130_fd_sc_hd__nand2_1 _23507_ (.A(_06829_),
    .B(_04257_),
    .Y(_06974_));
 sky130_fd_sc_hd__a21bo_1 _23508_ (.A1(_06974_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_06975_));
 sky130_fd_sc_hd__clkbuf_8 _23509_ (.A(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__mux2_1 _23510_ (.A0(_06530_),
    .A1(net2627),
    .S(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__clkbuf_1 _23511_ (.A(_06977_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _23512_ (.A0(_06538_),
    .A1(net2540),
    .S(_06976_),
    .X(_06978_));
 sky130_fd_sc_hd__clkbuf_1 _23513_ (.A(_06978_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _23514_ (.A0(_06540_),
    .A1(net2233),
    .S(_06976_),
    .X(_06979_));
 sky130_fd_sc_hd__clkbuf_1 _23515_ (.A(_06979_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _23516_ (.A0(_06542_),
    .A1(net2335),
    .S(_06976_),
    .X(_06980_));
 sky130_fd_sc_hd__clkbuf_1 _23517_ (.A(_06980_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _23518_ (.A0(_06544_),
    .A1(net2514),
    .S(_06976_),
    .X(_06981_));
 sky130_fd_sc_hd__clkbuf_1 _23519_ (.A(_06981_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _23520_ (.A0(_06546_),
    .A1(net2226),
    .S(_06976_),
    .X(_06982_));
 sky130_fd_sc_hd__clkbuf_1 _23521_ (.A(_06982_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _23522_ (.A0(_06548_),
    .A1(net2214),
    .S(_06976_),
    .X(_06983_));
 sky130_fd_sc_hd__clkbuf_1 _23523_ (.A(_06983_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _23524_ (.A0(_06550_),
    .A1(net3323),
    .S(_06976_),
    .X(_06984_));
 sky130_fd_sc_hd__clkbuf_1 _23525_ (.A(_06984_),
    .X(_01914_));
 sky130_fd_sc_hd__buf_4 _23526_ (.A(_06974_),
    .X(_06985_));
 sky130_fd_sc_hd__buf_4 _23527_ (.A(_06885_),
    .X(_06986_));
 sky130_fd_sc_hd__buf_4 _23528_ (.A(_06974_),
    .X(_06987_));
 sky130_fd_sc_hd__nand2_1 _23529_ (.A(_06987_),
    .B(_05010_),
    .Y(_06988_));
 sky130_fd_sc_hd__o211a_1 _23530_ (.A1(_05095_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__mux2_1 _23531_ (.A0(_06989_),
    .A1(net2599),
    .S(_06976_),
    .X(_06990_));
 sky130_fd_sc_hd__clkbuf_1 _23532_ (.A(_06990_),
    .X(_01915_));
 sky130_fd_sc_hd__nand2_1 _23533_ (.A(_06987_),
    .B(_05014_),
    .Y(_06991_));
 sky130_fd_sc_hd__o211a_1 _23534_ (.A1(_05101_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__mux2_1 _23535_ (.A0(_06992_),
    .A1(net2275),
    .S(_06976_),
    .X(_06993_));
 sky130_fd_sc_hd__clkbuf_1 _23536_ (.A(_06993_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _23537_ (.A(_06987_),
    .B(_05018_),
    .Y(_06994_));
 sky130_fd_sc_hd__o211a_1 _23538_ (.A1(_05105_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__mux2_1 _23539_ (.A0(_06995_),
    .A1(net2188),
    .S(_06976_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_1 _23540_ (.A(_06996_),
    .X(_01917_));
 sky130_fd_sc_hd__nand2_1 _23541_ (.A(_06987_),
    .B(_05022_),
    .Y(_06997_));
 sky130_fd_sc_hd__o211a_1 _23542_ (.A1(_05109_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__mux2_1 _23543_ (.A0(_06998_),
    .A1(net2457),
    .S(_06976_),
    .X(_06999_));
 sky130_fd_sc_hd__clkbuf_1 _23544_ (.A(_06999_),
    .X(_01918_));
 sky130_fd_sc_hd__nand2_1 _23545_ (.A(_06987_),
    .B(_05026_),
    .Y(_07000_));
 sky130_fd_sc_hd__o211a_1 _23546_ (.A1(_05113_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__mux2_1 _23547_ (.A0(_07001_),
    .A1(net2947),
    .S(_06976_),
    .X(_07002_));
 sky130_fd_sc_hd__clkbuf_1 _23548_ (.A(_07002_),
    .X(_01919_));
 sky130_fd_sc_hd__nand2_1 _23549_ (.A(_06987_),
    .B(_05030_),
    .Y(_07003_));
 sky130_fd_sc_hd__o211a_1 _23550_ (.A1(_05117_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__mux2_1 _23551_ (.A0(_07004_),
    .A1(net3189),
    .S(_06976_),
    .X(_07005_));
 sky130_fd_sc_hd__clkbuf_1 _23552_ (.A(_07005_),
    .X(_01920_));
 sky130_fd_sc_hd__nand2_1 _23553_ (.A(_06987_),
    .B(_05034_),
    .Y(_07006_));
 sky130_fd_sc_hd__o211a_1 _23554_ (.A1(_05121_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__mux2_1 _23555_ (.A0(_07007_),
    .A1(net3440),
    .S(_06976_),
    .X(_07008_));
 sky130_fd_sc_hd__clkbuf_1 _23556_ (.A(_07008_),
    .X(_01921_));
 sky130_fd_sc_hd__nand2_1 _23557_ (.A(_06987_),
    .B(_05038_),
    .Y(_07009_));
 sky130_fd_sc_hd__o211a_1 _23558_ (.A1(_05125_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__mux2_1 _23559_ (.A0(_07010_),
    .A1(net3594),
    .S(_06976_),
    .X(_07011_));
 sky130_fd_sc_hd__clkbuf_1 _23560_ (.A(_07011_),
    .X(_01922_));
 sky130_fd_sc_hd__o211a_1 _23561_ (.A1(_05129_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06988_),
    .X(_07012_));
 sky130_fd_sc_hd__clkbuf_8 _23562_ (.A(_06975_),
    .X(_07013_));
 sky130_fd_sc_hd__mux2_1 _23563_ (.A0(_07012_),
    .A1(net3358),
    .S(_07013_),
    .X(_07014_));
 sky130_fd_sc_hd__clkbuf_1 _23564_ (.A(_07014_),
    .X(_01923_));
 sky130_fd_sc_hd__o211a_1 _23565_ (.A1(_05134_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06991_),
    .X(_07015_));
 sky130_fd_sc_hd__mux2_1 _23566_ (.A0(_07015_),
    .A1(net2432),
    .S(_07013_),
    .X(_07016_));
 sky130_fd_sc_hd__clkbuf_1 _23567_ (.A(_07016_),
    .X(_01924_));
 sky130_fd_sc_hd__o211a_1 _23568_ (.A1(_05137_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06994_),
    .X(_07017_));
 sky130_fd_sc_hd__mux2_1 _23569_ (.A0(_07017_),
    .A1(net3377),
    .S(_07013_),
    .X(_07018_));
 sky130_fd_sc_hd__clkbuf_1 _23570_ (.A(_07018_),
    .X(_01925_));
 sky130_fd_sc_hd__o211a_1 _23571_ (.A1(_05140_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_06997_),
    .X(_07019_));
 sky130_fd_sc_hd__mux2_1 _23572_ (.A0(_07019_),
    .A1(net2436),
    .S(_07013_),
    .X(_07020_));
 sky130_fd_sc_hd__clkbuf_1 _23573_ (.A(_07020_),
    .X(_01926_));
 sky130_fd_sc_hd__o211a_1 _23574_ (.A1(_05143_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07000_),
    .X(_07021_));
 sky130_fd_sc_hd__mux2_1 _23575_ (.A0(_07021_),
    .A1(net2568),
    .S(_07013_),
    .X(_07022_));
 sky130_fd_sc_hd__clkbuf_1 _23576_ (.A(_07022_),
    .X(_01927_));
 sky130_fd_sc_hd__o211a_1 _23577_ (.A1(_05146_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07003_),
    .X(_07023_));
 sky130_fd_sc_hd__mux2_1 _23578_ (.A0(_07023_),
    .A1(net3590),
    .S(_07013_),
    .X(_07024_));
 sky130_fd_sc_hd__clkbuf_1 _23579_ (.A(_07024_),
    .X(_01928_));
 sky130_fd_sc_hd__o211a_1 _23580_ (.A1(_05149_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07006_),
    .X(_07025_));
 sky130_fd_sc_hd__mux2_1 _23581_ (.A0(_07025_),
    .A1(net3755),
    .S(_07013_),
    .X(_07026_));
 sky130_fd_sc_hd__clkbuf_1 _23582_ (.A(_07026_),
    .X(_01929_));
 sky130_fd_sc_hd__o211a_1 _23583_ (.A1(_05152_),
    .A2(_06985_),
    .B1(_06986_),
    .C1(_07009_),
    .X(_07027_));
 sky130_fd_sc_hd__mux2_1 _23584_ (.A0(_07027_),
    .A1(net2638),
    .S(_07013_),
    .X(_07028_));
 sky130_fd_sc_hd__clkbuf_1 _23585_ (.A(_07028_),
    .X(_01930_));
 sky130_fd_sc_hd__buf_4 _23586_ (.A(_06885_),
    .X(_07029_));
 sky130_fd_sc_hd__o211a_1 _23587_ (.A1(_05059_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_06988_),
    .X(_07030_));
 sky130_fd_sc_hd__mux2_1 _23588_ (.A0(_07030_),
    .A1(net3458),
    .S(_07013_),
    .X(_07031_));
 sky130_fd_sc_hd__clkbuf_1 _23589_ (.A(_07031_),
    .X(_01931_));
 sky130_fd_sc_hd__o211a_1 _23590_ (.A1(_05063_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_06991_),
    .X(_07032_));
 sky130_fd_sc_hd__mux2_1 _23591_ (.A0(_07032_),
    .A1(net3538),
    .S(_07013_),
    .X(_07033_));
 sky130_fd_sc_hd__clkbuf_1 _23592_ (.A(_07033_),
    .X(_01932_));
 sky130_fd_sc_hd__o211a_1 _23593_ (.A1(_05066_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_06994_),
    .X(_07034_));
 sky130_fd_sc_hd__mux2_1 _23594_ (.A0(_07034_),
    .A1(net3341),
    .S(_07013_),
    .X(_07035_));
 sky130_fd_sc_hd__clkbuf_1 _23595_ (.A(_07035_),
    .X(_01933_));
 sky130_fd_sc_hd__o211a_1 _23596_ (.A1(_05069_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_06997_),
    .X(_07036_));
 sky130_fd_sc_hd__mux2_1 _23597_ (.A0(_07036_),
    .A1(net3432),
    .S(_07013_),
    .X(_07037_));
 sky130_fd_sc_hd__clkbuf_1 _23598_ (.A(_07037_),
    .X(_01934_));
 sky130_fd_sc_hd__o211a_1 _23599_ (.A1(_05072_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_07000_),
    .X(_07038_));
 sky130_fd_sc_hd__mux2_1 _23600_ (.A0(_07038_),
    .A1(net3235),
    .S(_07013_),
    .X(_07039_));
 sky130_fd_sc_hd__clkbuf_1 _23601_ (.A(_07039_),
    .X(_01935_));
 sky130_fd_sc_hd__o211a_1 _23602_ (.A1(_05075_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_07003_),
    .X(_07040_));
 sky130_fd_sc_hd__mux2_1 _23603_ (.A0(_07040_),
    .A1(net3114),
    .S(_07013_),
    .X(_07041_));
 sky130_fd_sc_hd__clkbuf_1 _23604_ (.A(_07041_),
    .X(_01936_));
 sky130_fd_sc_hd__o211a_1 _23605_ (.A1(_05078_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_07006_),
    .X(_07042_));
 sky130_fd_sc_hd__mux2_1 _23606_ (.A0(_07042_),
    .A1(net3414),
    .S(_07013_),
    .X(_07043_));
 sky130_fd_sc_hd__clkbuf_1 _23607_ (.A(_07043_),
    .X(_01937_));
 sky130_fd_sc_hd__o211a_1 _23608_ (.A1(_05081_),
    .A2(_06987_),
    .B1(_07029_),
    .C1(_07009_),
    .X(_07044_));
 sky130_fd_sc_hd__mux2_1 _23609_ (.A0(_07044_),
    .A1(net3648),
    .S(_07013_),
    .X(_07045_));
 sky130_fd_sc_hd__clkbuf_1 _23610_ (.A(_07045_),
    .X(_01938_));
 sky130_fd_sc_hd__nand2_1 _23611_ (.A(_06829_),
    .B(_04333_),
    .Y(_07046_));
 sky130_fd_sc_hd__inv_2 _23612_ (.A(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__o21ai_4 _23613_ (.A1(_06755_),
    .A2(_07047_),
    .B1(_06020_),
    .Y(_07048_));
 sky130_fd_sc_hd__mux2_1 _23614_ (.A0(_06530_),
    .A1(net2831),
    .S(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__clkbuf_1 _23615_ (.A(_07049_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _23616_ (.A0(_06538_),
    .A1(net3006),
    .S(_07048_),
    .X(_07050_));
 sky130_fd_sc_hd__clkbuf_1 _23617_ (.A(_07050_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _23618_ (.A0(_06540_),
    .A1(net3737),
    .S(_07048_),
    .X(_07051_));
 sky130_fd_sc_hd__clkbuf_1 _23619_ (.A(_07051_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _23620_ (.A0(_06542_),
    .A1(net3316),
    .S(_07048_),
    .X(_07052_));
 sky130_fd_sc_hd__clkbuf_1 _23621_ (.A(_07052_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _23622_ (.A0(_06544_),
    .A1(net2559),
    .S(_07048_),
    .X(_07053_));
 sky130_fd_sc_hd__clkbuf_1 _23623_ (.A(_07053_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _23624_ (.A0(_06546_),
    .A1(net2592),
    .S(_07048_),
    .X(_07054_));
 sky130_fd_sc_hd__clkbuf_1 _23625_ (.A(_07054_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _23626_ (.A0(_06548_),
    .A1(net3239),
    .S(_07048_),
    .X(_07055_));
 sky130_fd_sc_hd__clkbuf_1 _23627_ (.A(_07055_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _23628_ (.A0(_06550_),
    .A1(net2120),
    .S(_07048_),
    .X(_07056_));
 sky130_fd_sc_hd__clkbuf_1 _23629_ (.A(_07056_),
    .X(_01946_));
 sky130_fd_sc_hd__buf_4 _23630_ (.A(_07048_),
    .X(_07057_));
 sky130_fd_sc_hd__buf_4 _23631_ (.A(_07047_),
    .X(_07058_));
 sky130_fd_sc_hd__buf_4 _23632_ (.A(_07047_),
    .X(_07059_));
 sky130_fd_sc_hd__nor2_1 _23633_ (.A(_05583_),
    .B(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__a211o_1 _23634_ (.A1(_05484_),
    .A2(_07058_),
    .B1(_06800_),
    .C1(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__buf_4 _23635_ (.A(_07048_),
    .X(_07062_));
 sky130_fd_sc_hd__nand2_1 _23636_ (.A(_07062_),
    .B(net812),
    .Y(_07063_));
 sky130_fd_sc_hd__o21ai_1 _23637_ (.A1(_07057_),
    .A2(_07061_),
    .B1(net813),
    .Y(_01947_));
 sky130_fd_sc_hd__nor2_1 _23638_ (.A(_05589_),
    .B(_07059_),
    .Y(_07064_));
 sky130_fd_sc_hd__a211o_1 _23639_ (.A1(_05491_),
    .A2(_07058_),
    .B1(_06800_),
    .C1(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__nand2_1 _23640_ (.A(_07062_),
    .B(net1592),
    .Y(_07066_));
 sky130_fd_sc_hd__o21ai_1 _23641_ (.A1(_07057_),
    .A2(_07065_),
    .B1(net1593),
    .Y(_01948_));
 sky130_fd_sc_hd__buf_4 _23642_ (.A(_05892_),
    .X(_07067_));
 sky130_fd_sc_hd__nor2_1 _23643_ (.A(_05593_),
    .B(_07059_),
    .Y(_07068_));
 sky130_fd_sc_hd__a211o_1 _23644_ (.A1(_05495_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__nand2_1 _23645_ (.A(_07062_),
    .B(net1472),
    .Y(_07070_));
 sky130_fd_sc_hd__o21ai_1 _23646_ (.A1(_07057_),
    .A2(_07069_),
    .B1(net1473),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_1 _23647_ (.A(_05597_),
    .B(_07059_),
    .Y(_07071_));
 sky130_fd_sc_hd__a211o_1 _23648_ (.A1(_05500_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07071_),
    .X(_07072_));
 sky130_fd_sc_hd__nand2_1 _23649_ (.A(_07062_),
    .B(net1772),
    .Y(_07073_));
 sky130_fd_sc_hd__o21ai_1 _23650_ (.A1(_07057_),
    .A2(_07072_),
    .B1(net1773),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_1 _23651_ (.A(_05601_),
    .B(_07059_),
    .Y(_07074_));
 sky130_fd_sc_hd__a211o_1 _23652_ (.A1(_05504_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__nand2_1 _23653_ (.A(_07062_),
    .B(net1798),
    .Y(_07076_));
 sky130_fd_sc_hd__o21ai_1 _23654_ (.A1(_07057_),
    .A2(_07075_),
    .B1(net1799),
    .Y(_01951_));
 sky130_fd_sc_hd__nor2_1 _23655_ (.A(_05605_),
    .B(_07059_),
    .Y(_07077_));
 sky130_fd_sc_hd__a211o_1 _23656_ (.A1(_05508_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07077_),
    .X(_07078_));
 sky130_fd_sc_hd__nand2_1 _23657_ (.A(_07062_),
    .B(net1146),
    .Y(_07079_));
 sky130_fd_sc_hd__o21ai_1 _23658_ (.A1(_07057_),
    .A2(_07078_),
    .B1(net1147),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _23659_ (.A(_05609_),
    .B(_07059_),
    .Y(_07080_));
 sky130_fd_sc_hd__a211o_1 _23660_ (.A1(_05512_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__nand2_1 _23661_ (.A(_07062_),
    .B(net1796),
    .Y(_07082_));
 sky130_fd_sc_hd__o21ai_1 _23662_ (.A1(_07057_),
    .A2(_07081_),
    .B1(net1797),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _23663_ (.A(_05613_),
    .B(_07059_),
    .Y(_07083_));
 sky130_fd_sc_hd__a211o_1 _23664_ (.A1(_05516_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__nand2_1 _23665_ (.A(_07062_),
    .B(net1923),
    .Y(_07085_));
 sky130_fd_sc_hd__o21ai_1 _23666_ (.A1(_07057_),
    .A2(_07084_),
    .B1(net1924),
    .Y(_01954_));
 sky130_fd_sc_hd__buf_4 _23667_ (.A(_07048_),
    .X(_07086_));
 sky130_fd_sc_hd__a211o_1 _23668_ (.A1(_05521_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07060_),
    .X(_07087_));
 sky130_fd_sc_hd__nand2_1 _23669_ (.A(_07062_),
    .B(net1666),
    .Y(_07088_));
 sky130_fd_sc_hd__o21ai_1 _23670_ (.A1(_07086_),
    .A2(_07087_),
    .B1(net1667),
    .Y(_01955_));
 sky130_fd_sc_hd__a211o_1 _23671_ (.A1(_05524_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07064_),
    .X(_07089_));
 sky130_fd_sc_hd__nand2_1 _23672_ (.A(_07062_),
    .B(net1794),
    .Y(_07090_));
 sky130_fd_sc_hd__o21ai_1 _23673_ (.A1(_07086_),
    .A2(_07089_),
    .B1(net1795),
    .Y(_01956_));
 sky130_fd_sc_hd__a211o_1 _23674_ (.A1(_05527_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07068_),
    .X(_07091_));
 sky130_fd_sc_hd__nand2_1 _23675_ (.A(_07062_),
    .B(net1496),
    .Y(_07092_));
 sky130_fd_sc_hd__o21ai_1 _23676_ (.A1(_07086_),
    .A2(_07091_),
    .B1(net1497),
    .Y(_01957_));
 sky130_fd_sc_hd__a211o_1 _23677_ (.A1(_05530_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07071_),
    .X(_07093_));
 sky130_fd_sc_hd__nand2_1 _23678_ (.A(_07062_),
    .B(net1948),
    .Y(_07094_));
 sky130_fd_sc_hd__o21ai_1 _23679_ (.A1(_07086_),
    .A2(_07093_),
    .B1(net1949),
    .Y(_01958_));
 sky130_fd_sc_hd__a211o_1 _23680_ (.A1(_05533_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07074_),
    .X(_07095_));
 sky130_fd_sc_hd__nand2_1 _23681_ (.A(_07062_),
    .B(net1931),
    .Y(_07096_));
 sky130_fd_sc_hd__o21ai_1 _23682_ (.A1(_07086_),
    .A2(_07095_),
    .B1(_07096_),
    .Y(_01959_));
 sky130_fd_sc_hd__a211o_1 _23683_ (.A1(_05536_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07077_),
    .X(_07097_));
 sky130_fd_sc_hd__nand2_1 _23684_ (.A(_07062_),
    .B(net1432),
    .Y(_07098_));
 sky130_fd_sc_hd__o21ai_1 _23685_ (.A1(_07086_),
    .A2(_07097_),
    .B1(net1433),
    .Y(_01960_));
 sky130_fd_sc_hd__a211o_1 _23686_ (.A1(_05539_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07080_),
    .X(_07099_));
 sky130_fd_sc_hd__nand2_1 _23687_ (.A(_07062_),
    .B(net1820),
    .Y(_07100_));
 sky130_fd_sc_hd__o21ai_1 _23688_ (.A1(_07086_),
    .A2(_07099_),
    .B1(net1821),
    .Y(_01961_));
 sky130_fd_sc_hd__a211o_1 _23689_ (.A1(_05542_),
    .A2(_07058_),
    .B1(_07067_),
    .C1(_07083_),
    .X(_07101_));
 sky130_fd_sc_hd__nand2_1 _23690_ (.A(_07062_),
    .B(net1972),
    .Y(_07102_));
 sky130_fd_sc_hd__o21ai_1 _23691_ (.A1(_07086_),
    .A2(_07101_),
    .B1(_07102_),
    .Y(_01962_));
 sky130_fd_sc_hd__a211o_1 _23692_ (.A1(_05545_),
    .A2(_07059_),
    .B1(_07067_),
    .C1(_07060_),
    .X(_07103_));
 sky130_fd_sc_hd__nand2_1 _23693_ (.A(_07057_),
    .B(net554),
    .Y(_07104_));
 sky130_fd_sc_hd__o21ai_1 _23694_ (.A1(_07086_),
    .A2(_07103_),
    .B1(net555),
    .Y(_01963_));
 sky130_fd_sc_hd__a211o_1 _23695_ (.A1(_05548_),
    .A2(_07059_),
    .B1(_07067_),
    .C1(_07064_),
    .X(_07105_));
 sky130_fd_sc_hd__nand2_1 _23696_ (.A(_07057_),
    .B(net392),
    .Y(_07106_));
 sky130_fd_sc_hd__o21ai_1 _23697_ (.A1(_07086_),
    .A2(_07105_),
    .B1(net393),
    .Y(_01964_));
 sky130_fd_sc_hd__clkbuf_8 _23698_ (.A(_05892_),
    .X(_07107_));
 sky130_fd_sc_hd__a211o_1 _23699_ (.A1(_05551_),
    .A2(_07059_),
    .B1(_07107_),
    .C1(_07068_),
    .X(_07108_));
 sky130_fd_sc_hd__nand2_1 _23700_ (.A(_07057_),
    .B(net1050),
    .Y(_07109_));
 sky130_fd_sc_hd__o21ai_1 _23701_ (.A1(_07086_),
    .A2(_07108_),
    .B1(net1051),
    .Y(_01965_));
 sky130_fd_sc_hd__a211o_1 _23702_ (.A1(_05555_),
    .A2(_07059_),
    .B1(_07107_),
    .C1(_07071_),
    .X(_07110_));
 sky130_fd_sc_hd__nand2_1 _23703_ (.A(_07057_),
    .B(net1376),
    .Y(_07111_));
 sky130_fd_sc_hd__o21ai_1 _23704_ (.A1(_07086_),
    .A2(_07110_),
    .B1(net1377),
    .Y(_01966_));
 sky130_fd_sc_hd__a211o_1 _23705_ (.A1(_05558_),
    .A2(_07059_),
    .B1(_07107_),
    .C1(_07074_),
    .X(_07112_));
 sky130_fd_sc_hd__nand2_1 _23706_ (.A(_07057_),
    .B(net1616),
    .Y(_07113_));
 sky130_fd_sc_hd__o21ai_1 _23707_ (.A1(_07086_),
    .A2(_07112_),
    .B1(net1617),
    .Y(_01967_));
 sky130_fd_sc_hd__a211o_1 _23708_ (.A1(_05561_),
    .A2(_07059_),
    .B1(_07107_),
    .C1(_07077_),
    .X(_07114_));
 sky130_fd_sc_hd__nand2_1 _23709_ (.A(_07057_),
    .B(net1860),
    .Y(_07115_));
 sky130_fd_sc_hd__o21ai_1 _23710_ (.A1(_07086_),
    .A2(_07114_),
    .B1(net1861),
    .Y(_01968_));
 sky130_fd_sc_hd__a211o_1 _23711_ (.A1(_05564_),
    .A2(_07059_),
    .B1(_07107_),
    .C1(_07080_),
    .X(_07116_));
 sky130_fd_sc_hd__nand2_1 _23712_ (.A(_07057_),
    .B(net1978),
    .Y(_07117_));
 sky130_fd_sc_hd__o21ai_1 _23713_ (.A1(_07086_),
    .A2(_07116_),
    .B1(_07117_),
    .Y(_01969_));
 sky130_fd_sc_hd__a211o_1 _23714_ (.A1(_05567_),
    .A2(_07059_),
    .B1(_07107_),
    .C1(_07083_),
    .X(_07118_));
 sky130_fd_sc_hd__nand2_1 _23715_ (.A(_07057_),
    .B(net1977),
    .Y(_07119_));
 sky130_fd_sc_hd__o21ai_1 _23716_ (.A1(_07086_),
    .A2(_07118_),
    .B1(_07119_),
    .Y(_01970_));
 sky130_fd_sc_hd__and2_2 _23717_ (.A(_03516_),
    .B(_06531_),
    .X(_07120_));
 sky130_fd_sc_hd__nand2_1 _23718_ (.A(_07120_),
    .B(_04104_),
    .Y(_07121_));
 sky130_fd_sc_hd__a21bo_1 _23719_ (.A1(_07121_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_07122_));
 sky130_fd_sc_hd__clkbuf_8 _23720_ (.A(_07122_),
    .X(_07123_));
 sky130_fd_sc_hd__mux2_1 _23721_ (.A0(_06530_),
    .A1(net3272),
    .S(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__clkbuf_1 _23722_ (.A(_07124_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _23723_ (.A0(_06538_),
    .A1(net2182),
    .S(_07123_),
    .X(_07125_));
 sky130_fd_sc_hd__clkbuf_1 _23724_ (.A(_07125_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _23725_ (.A0(_06540_),
    .A1(net3439),
    .S(_07123_),
    .X(_07126_));
 sky130_fd_sc_hd__clkbuf_1 _23726_ (.A(_07126_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _23727_ (.A0(_06542_),
    .A1(net2045),
    .S(_07123_),
    .X(_07127_));
 sky130_fd_sc_hd__clkbuf_1 _23728_ (.A(_07127_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _23729_ (.A0(_06544_),
    .A1(net2023),
    .S(_07123_),
    .X(_07128_));
 sky130_fd_sc_hd__clkbuf_1 _23730_ (.A(_07128_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _23731_ (.A0(_06546_),
    .A1(net2089),
    .S(_07123_),
    .X(_07129_));
 sky130_fd_sc_hd__clkbuf_1 _23732_ (.A(_07129_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _23733_ (.A0(_06548_),
    .A1(net2122),
    .S(_07123_),
    .X(_07130_));
 sky130_fd_sc_hd__clkbuf_1 _23734_ (.A(_07130_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _23735_ (.A0(_06550_),
    .A1(net2309),
    .S(_07123_),
    .X(_07131_));
 sky130_fd_sc_hd__clkbuf_1 _23736_ (.A(_07131_),
    .X(_01978_));
 sky130_fd_sc_hd__buf_4 _23737_ (.A(_07121_),
    .X(_07132_));
 sky130_fd_sc_hd__buf_4 _23738_ (.A(_07121_),
    .X(_07133_));
 sky130_fd_sc_hd__nand2_1 _23739_ (.A(_07133_),
    .B(_05010_),
    .Y(_07134_));
 sky130_fd_sc_hd__o211a_1 _23740_ (.A1(_05095_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__mux2_1 _23741_ (.A0(_07135_),
    .A1(net2902),
    .S(_07123_),
    .X(_07136_));
 sky130_fd_sc_hd__clkbuf_1 _23742_ (.A(_07136_),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_1 _23743_ (.A(_07133_),
    .B(_05014_),
    .Y(_07137_));
 sky130_fd_sc_hd__o211a_1 _23744_ (.A1(_05101_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__mux2_1 _23745_ (.A0(_07138_),
    .A1(net2096),
    .S(_07123_),
    .X(_07139_));
 sky130_fd_sc_hd__clkbuf_1 _23746_ (.A(_07139_),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_1 _23747_ (.A(_07133_),
    .B(_05018_),
    .Y(_07140_));
 sky130_fd_sc_hd__o211a_1 _23748_ (.A1(_05105_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__mux2_1 _23749_ (.A0(_07141_),
    .A1(net2756),
    .S(_07123_),
    .X(_07142_));
 sky130_fd_sc_hd__clkbuf_1 _23750_ (.A(_07142_),
    .X(_01981_));
 sky130_fd_sc_hd__nand2_1 _23751_ (.A(_07133_),
    .B(_05022_),
    .Y(_07143_));
 sky130_fd_sc_hd__o211a_1 _23752_ (.A1(_05109_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__mux2_1 _23753_ (.A0(_07144_),
    .A1(net2060),
    .S(_07123_),
    .X(_07145_));
 sky130_fd_sc_hd__clkbuf_1 _23754_ (.A(_07145_),
    .X(_01982_));
 sky130_fd_sc_hd__nand2_1 _23755_ (.A(_07133_),
    .B(_05026_),
    .Y(_07146_));
 sky130_fd_sc_hd__o211a_1 _23756_ (.A1(_05113_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__mux2_1 _23757_ (.A0(_07147_),
    .A1(net2054),
    .S(_07123_),
    .X(_07148_));
 sky130_fd_sc_hd__clkbuf_1 _23758_ (.A(_07148_),
    .X(_01983_));
 sky130_fd_sc_hd__nand2_1 _23759_ (.A(_07133_),
    .B(_05030_),
    .Y(_07149_));
 sky130_fd_sc_hd__o211a_1 _23760_ (.A1(_05117_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__mux2_1 _23761_ (.A0(_07150_),
    .A1(net2193),
    .S(_07123_),
    .X(_07151_));
 sky130_fd_sc_hd__clkbuf_1 _23762_ (.A(_07151_),
    .X(_01984_));
 sky130_fd_sc_hd__nand2_1 _23763_ (.A(_07133_),
    .B(_05034_),
    .Y(_07152_));
 sky130_fd_sc_hd__o211a_1 _23764_ (.A1(_05121_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__mux2_1 _23765_ (.A0(_07153_),
    .A1(net2220),
    .S(_07123_),
    .X(_07154_));
 sky130_fd_sc_hd__clkbuf_1 _23766_ (.A(_07154_),
    .X(_01985_));
 sky130_fd_sc_hd__nand2_1 _23767_ (.A(_07133_),
    .B(_05038_),
    .Y(_07155_));
 sky130_fd_sc_hd__o211a_1 _23768_ (.A1(_05125_),
    .A2(_07132_),
    .B1(_07029_),
    .C1(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__mux2_1 _23769_ (.A0(_07156_),
    .A1(net2077),
    .S(_07123_),
    .X(_07157_));
 sky130_fd_sc_hd__clkbuf_1 _23770_ (.A(_07157_),
    .X(_01986_));
 sky130_fd_sc_hd__buf_4 _23771_ (.A(_06885_),
    .X(_07158_));
 sky130_fd_sc_hd__o211a_1 _23772_ (.A1(_05129_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07134_),
    .X(_07159_));
 sky130_fd_sc_hd__clkbuf_8 _23773_ (.A(_07122_),
    .X(_07160_));
 sky130_fd_sc_hd__mux2_1 _23774_ (.A0(_07159_),
    .A1(net2132),
    .S(_07160_),
    .X(_07161_));
 sky130_fd_sc_hd__clkbuf_1 _23775_ (.A(_07161_),
    .X(_01987_));
 sky130_fd_sc_hd__o211a_1 _23776_ (.A1(_05134_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07137_),
    .X(_07162_));
 sky130_fd_sc_hd__mux2_1 _23777_ (.A0(_07162_),
    .A1(net2090),
    .S(_07160_),
    .X(_07163_));
 sky130_fd_sc_hd__clkbuf_1 _23778_ (.A(_07163_),
    .X(_01988_));
 sky130_fd_sc_hd__o211a_1 _23779_ (.A1(_05137_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07140_),
    .X(_07164_));
 sky130_fd_sc_hd__mux2_1 _23780_ (.A0(_07164_),
    .A1(net2043),
    .S(_07160_),
    .X(_07165_));
 sky130_fd_sc_hd__clkbuf_1 _23781_ (.A(_07165_),
    .X(_01989_));
 sky130_fd_sc_hd__o211a_1 _23782_ (.A1(_05140_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07143_),
    .X(_07166_));
 sky130_fd_sc_hd__mux2_1 _23783_ (.A0(_07166_),
    .A1(net2164),
    .S(_07160_),
    .X(_07167_));
 sky130_fd_sc_hd__clkbuf_1 _23784_ (.A(_07167_),
    .X(_01990_));
 sky130_fd_sc_hd__o211a_1 _23785_ (.A1(_05143_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07146_),
    .X(_07168_));
 sky130_fd_sc_hd__mux2_1 _23786_ (.A0(_07168_),
    .A1(net2266),
    .S(_07160_),
    .X(_07169_));
 sky130_fd_sc_hd__clkbuf_1 _23787_ (.A(_07169_),
    .X(_01991_));
 sky130_fd_sc_hd__o211a_1 _23788_ (.A1(_05146_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07149_),
    .X(_07170_));
 sky130_fd_sc_hd__mux2_1 _23789_ (.A0(_07170_),
    .A1(net2127),
    .S(_07160_),
    .X(_07171_));
 sky130_fd_sc_hd__clkbuf_1 _23790_ (.A(_07171_),
    .X(_01992_));
 sky130_fd_sc_hd__o211a_1 _23791_ (.A1(_05149_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07152_),
    .X(_07172_));
 sky130_fd_sc_hd__mux2_1 _23792_ (.A0(_07172_),
    .A1(net2115),
    .S(_07160_),
    .X(_07173_));
 sky130_fd_sc_hd__clkbuf_1 _23793_ (.A(_07173_),
    .X(_01993_));
 sky130_fd_sc_hd__o211a_1 _23794_ (.A1(_05152_),
    .A2(_07132_),
    .B1(_07158_),
    .C1(_07155_),
    .X(_07174_));
 sky130_fd_sc_hd__mux2_1 _23795_ (.A0(_07174_),
    .A1(net2191),
    .S(_07160_),
    .X(_07175_));
 sky130_fd_sc_hd__clkbuf_1 _23796_ (.A(_07175_),
    .X(_01994_));
 sky130_fd_sc_hd__o211a_1 _23797_ (.A1(_05059_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07134_),
    .X(_07176_));
 sky130_fd_sc_hd__mux2_1 _23798_ (.A0(_07176_),
    .A1(net2142),
    .S(_07160_),
    .X(_07177_));
 sky130_fd_sc_hd__clkbuf_1 _23799_ (.A(_07177_),
    .X(_01995_));
 sky130_fd_sc_hd__o211a_1 _23800_ (.A1(_05063_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07137_),
    .X(_07178_));
 sky130_fd_sc_hd__mux2_1 _23801_ (.A0(_07178_),
    .A1(net2140),
    .S(_07160_),
    .X(_07179_));
 sky130_fd_sc_hd__clkbuf_1 _23802_ (.A(_07179_),
    .X(_01996_));
 sky130_fd_sc_hd__o211a_1 _23803_ (.A1(_05066_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07140_),
    .X(_07180_));
 sky130_fd_sc_hd__mux2_1 _23804_ (.A0(_07180_),
    .A1(net2167),
    .S(_07160_),
    .X(_07181_));
 sky130_fd_sc_hd__clkbuf_1 _23805_ (.A(_07181_),
    .X(_01997_));
 sky130_fd_sc_hd__o211a_1 _23806_ (.A1(_05069_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07143_),
    .X(_07182_));
 sky130_fd_sc_hd__mux2_1 _23807_ (.A0(_07182_),
    .A1(net2165),
    .S(_07160_),
    .X(_07183_));
 sky130_fd_sc_hd__clkbuf_1 _23808_ (.A(_07183_),
    .X(_01998_));
 sky130_fd_sc_hd__o211a_1 _23809_ (.A1(_05072_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07146_),
    .X(_07184_));
 sky130_fd_sc_hd__mux2_1 _23810_ (.A0(_07184_),
    .A1(net2071),
    .S(_07160_),
    .X(_07185_));
 sky130_fd_sc_hd__clkbuf_1 _23811_ (.A(_07185_),
    .X(_01999_));
 sky130_fd_sc_hd__o211a_1 _23812_ (.A1(_05075_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07149_),
    .X(_07186_));
 sky130_fd_sc_hd__mux2_1 _23813_ (.A0(_07186_),
    .A1(net2072),
    .S(_07160_),
    .X(_07187_));
 sky130_fd_sc_hd__clkbuf_1 _23814_ (.A(_07187_),
    .X(_02000_));
 sky130_fd_sc_hd__o211a_1 _23815_ (.A1(_05078_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07152_),
    .X(_07188_));
 sky130_fd_sc_hd__mux2_1 _23816_ (.A0(_07188_),
    .A1(net2095),
    .S(_07160_),
    .X(_07189_));
 sky130_fd_sc_hd__clkbuf_1 _23817_ (.A(_07189_),
    .X(_02001_));
 sky130_fd_sc_hd__o211a_1 _23818_ (.A1(_05081_),
    .A2(_07133_),
    .B1(_07158_),
    .C1(_07155_),
    .X(_07190_));
 sky130_fd_sc_hd__mux2_1 _23819_ (.A0(_07190_),
    .A1(net2039),
    .S(_07160_),
    .X(_07191_));
 sky130_fd_sc_hd__clkbuf_1 _23820_ (.A(_07191_),
    .X(_02002_));
 sky130_fd_sc_hd__nand2_1 _23821_ (.A(_07120_),
    .B(_04183_),
    .Y(_07192_));
 sky130_fd_sc_hd__a21bo_1 _23822_ (.A1(_07192_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_07193_));
 sky130_fd_sc_hd__clkbuf_8 _23823_ (.A(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__mux2_1 _23824_ (.A0(_06530_),
    .A1(net2106),
    .S(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__clkbuf_1 _23825_ (.A(_07195_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _23826_ (.A0(_06538_),
    .A1(net2174),
    .S(_07194_),
    .X(_07196_));
 sky130_fd_sc_hd__clkbuf_1 _23827_ (.A(_07196_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _23828_ (.A0(_06540_),
    .A1(net2170),
    .S(_07194_),
    .X(_07197_));
 sky130_fd_sc_hd__clkbuf_1 _23829_ (.A(_07197_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _23830_ (.A0(_06542_),
    .A1(net2067),
    .S(_07194_),
    .X(_07198_));
 sky130_fd_sc_hd__clkbuf_1 _23831_ (.A(_07198_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _23832_ (.A0(_06544_),
    .A1(net2107),
    .S(_07194_),
    .X(_07199_));
 sky130_fd_sc_hd__clkbuf_1 _23833_ (.A(_07199_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _23834_ (.A0(_06546_),
    .A1(net3048),
    .S(_07194_),
    .X(_07200_));
 sky130_fd_sc_hd__clkbuf_1 _23835_ (.A(_07200_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _23836_ (.A0(_06548_),
    .A1(net2888),
    .S(_07194_),
    .X(_07201_));
 sky130_fd_sc_hd__clkbuf_1 _23837_ (.A(_07201_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _23838_ (.A0(_06550_),
    .A1(net2062),
    .S(_07194_),
    .X(_07202_));
 sky130_fd_sc_hd__clkbuf_1 _23839_ (.A(_07202_),
    .X(_02010_));
 sky130_fd_sc_hd__buf_4 _23840_ (.A(_07192_),
    .X(_07203_));
 sky130_fd_sc_hd__buf_4 _23841_ (.A(_06885_),
    .X(_07204_));
 sky130_fd_sc_hd__buf_4 _23842_ (.A(_07192_),
    .X(_07205_));
 sky130_fd_sc_hd__nand2_1 _23843_ (.A(_07205_),
    .B(_12184_),
    .Y(_07206_));
 sky130_fd_sc_hd__o211a_1 _23844_ (.A1(_05095_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07206_),
    .X(_07207_));
 sky130_fd_sc_hd__mux2_1 _23845_ (.A0(_07207_),
    .A1(net2271),
    .S(_07194_),
    .X(_07208_));
 sky130_fd_sc_hd__clkbuf_1 _23846_ (.A(_07208_),
    .X(_02011_));
 sky130_fd_sc_hd__nand2_1 _23847_ (.A(_07205_),
    .B(_12197_),
    .Y(_07209_));
 sky130_fd_sc_hd__o211a_1 _23848_ (.A1(_05101_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__mux2_1 _23849_ (.A0(_07210_),
    .A1(net2645),
    .S(_07194_),
    .X(_07211_));
 sky130_fd_sc_hd__clkbuf_1 _23850_ (.A(_07211_),
    .X(_02012_));
 sky130_fd_sc_hd__nand2_1 _23851_ (.A(_07205_),
    .B(_12205_),
    .Y(_07212_));
 sky130_fd_sc_hd__o211a_1 _23852_ (.A1(_05105_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__mux2_1 _23853_ (.A0(_07213_),
    .A1(net3375),
    .S(_07194_),
    .X(_07214_));
 sky130_fd_sc_hd__clkbuf_1 _23854_ (.A(_07214_),
    .X(_02013_));
 sky130_fd_sc_hd__nand2_1 _23855_ (.A(_07205_),
    .B(_12213_),
    .Y(_07215_));
 sky130_fd_sc_hd__o211a_1 _23856_ (.A1(_05109_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07215_),
    .X(_07216_));
 sky130_fd_sc_hd__mux2_1 _23857_ (.A0(_07216_),
    .A1(net2301),
    .S(_07194_),
    .X(_07217_));
 sky130_fd_sc_hd__clkbuf_1 _23858_ (.A(_07217_),
    .X(_02014_));
 sky130_fd_sc_hd__nand2_1 _23859_ (.A(_07205_),
    .B(_12221_),
    .Y(_07218_));
 sky130_fd_sc_hd__o211a_1 _23860_ (.A1(_05113_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__mux2_1 _23861_ (.A0(_07219_),
    .A1(net3220),
    .S(_07194_),
    .X(_07220_));
 sky130_fd_sc_hd__clkbuf_1 _23862_ (.A(_07220_),
    .X(_02015_));
 sky130_fd_sc_hd__nand2_1 _23863_ (.A(_07205_),
    .B(_12229_),
    .Y(_07221_));
 sky130_fd_sc_hd__o211a_1 _23864_ (.A1(_05117_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__mux2_1 _23865_ (.A0(_07222_),
    .A1(net2104),
    .S(_07194_),
    .X(_07223_));
 sky130_fd_sc_hd__clkbuf_1 _23866_ (.A(_07223_),
    .X(_02016_));
 sky130_fd_sc_hd__nand2_1 _23867_ (.A(_07205_),
    .B(_12237_),
    .Y(_07224_));
 sky130_fd_sc_hd__o211a_1 _23868_ (.A1(_05121_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__mux2_1 _23869_ (.A0(_07225_),
    .A1(net2066),
    .S(_07194_),
    .X(_07226_));
 sky130_fd_sc_hd__clkbuf_1 _23870_ (.A(_07226_),
    .X(_02017_));
 sky130_fd_sc_hd__nand2_1 _23871_ (.A(_07205_),
    .B(_12245_),
    .Y(_07227_));
 sky130_fd_sc_hd__o211a_1 _23872_ (.A1(_05125_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__mux2_1 _23873_ (.A0(_07228_),
    .A1(net2129),
    .S(_07194_),
    .X(_07229_));
 sky130_fd_sc_hd__clkbuf_1 _23874_ (.A(_07229_),
    .X(_02018_));
 sky130_fd_sc_hd__o211a_1 _23875_ (.A1(_05129_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07206_),
    .X(_07230_));
 sky130_fd_sc_hd__clkbuf_8 _23876_ (.A(_07193_),
    .X(_07231_));
 sky130_fd_sc_hd__mux2_1 _23877_ (.A0(_07230_),
    .A1(net3417),
    .S(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__clkbuf_1 _23878_ (.A(_07232_),
    .X(_02019_));
 sky130_fd_sc_hd__o211a_1 _23879_ (.A1(_05134_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07209_),
    .X(_07233_));
 sky130_fd_sc_hd__mux2_1 _23880_ (.A0(_07233_),
    .A1(net2399),
    .S(_07231_),
    .X(_07234_));
 sky130_fd_sc_hd__clkbuf_1 _23881_ (.A(_07234_),
    .X(_02020_));
 sky130_fd_sc_hd__o211a_1 _23882_ (.A1(_05137_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07212_),
    .X(_07235_));
 sky130_fd_sc_hd__mux2_1 _23883_ (.A0(_07235_),
    .A1(net3567),
    .S(_07231_),
    .X(_07236_));
 sky130_fd_sc_hd__clkbuf_1 _23884_ (.A(_07236_),
    .X(_02021_));
 sky130_fd_sc_hd__o211a_1 _23885_ (.A1(_05140_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07215_),
    .X(_07237_));
 sky130_fd_sc_hd__mux2_1 _23886_ (.A0(_07237_),
    .A1(net3634),
    .S(_07231_),
    .X(_07238_));
 sky130_fd_sc_hd__clkbuf_1 _23887_ (.A(_07238_),
    .X(_02022_));
 sky130_fd_sc_hd__o211a_1 _23888_ (.A1(_05143_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07218_),
    .X(_07239_));
 sky130_fd_sc_hd__mux2_1 _23889_ (.A0(_07239_),
    .A1(net3631),
    .S(_07231_),
    .X(_07240_));
 sky130_fd_sc_hd__clkbuf_1 _23890_ (.A(_07240_),
    .X(_02023_));
 sky130_fd_sc_hd__o211a_1 _23891_ (.A1(_05146_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07221_),
    .X(_07241_));
 sky130_fd_sc_hd__mux2_1 _23892_ (.A0(_07241_),
    .A1(net2482),
    .S(_07231_),
    .X(_07242_));
 sky130_fd_sc_hd__clkbuf_1 _23893_ (.A(_07242_),
    .X(_02024_));
 sky130_fd_sc_hd__o211a_1 _23894_ (.A1(_05149_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07224_),
    .X(_07243_));
 sky130_fd_sc_hd__mux2_1 _23895_ (.A0(_07243_),
    .A1(net2327),
    .S(_07231_),
    .X(_07244_));
 sky130_fd_sc_hd__clkbuf_1 _23896_ (.A(_07244_),
    .X(_02025_));
 sky130_fd_sc_hd__o211a_1 _23897_ (.A1(_05152_),
    .A2(_07203_),
    .B1(_07204_),
    .C1(_07227_),
    .X(_07245_));
 sky130_fd_sc_hd__mux2_1 _23898_ (.A0(_07245_),
    .A1(net2409),
    .S(_07231_),
    .X(_07246_));
 sky130_fd_sc_hd__clkbuf_1 _23899_ (.A(_07246_),
    .X(_02026_));
 sky130_fd_sc_hd__buf_4 _23900_ (.A(_06885_),
    .X(_07247_));
 sky130_fd_sc_hd__o211a_1 _23901_ (.A1(_12169_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07206_),
    .X(_07248_));
 sky130_fd_sc_hd__mux2_1 _23902_ (.A0(_07248_),
    .A1(net2442),
    .S(_07231_),
    .X(_07249_));
 sky130_fd_sc_hd__clkbuf_1 _23903_ (.A(_07249_),
    .X(_02027_));
 sky130_fd_sc_hd__o211a_1 _23904_ (.A1(_12194_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07209_),
    .X(_07250_));
 sky130_fd_sc_hd__mux2_1 _23905_ (.A0(_07250_),
    .A1(net3447),
    .S(_07231_),
    .X(_07251_));
 sky130_fd_sc_hd__clkbuf_1 _23906_ (.A(_07251_),
    .X(_02028_));
 sky130_fd_sc_hd__o211a_1 _23907_ (.A1(_12202_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07212_),
    .X(_07252_));
 sky130_fd_sc_hd__mux2_1 _23908_ (.A0(_07252_),
    .A1(net2647),
    .S(_07231_),
    .X(_07253_));
 sky130_fd_sc_hd__clkbuf_1 _23909_ (.A(_07253_),
    .X(_02029_));
 sky130_fd_sc_hd__o211a_1 _23910_ (.A1(_12210_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07215_),
    .X(_07254_));
 sky130_fd_sc_hd__mux2_1 _23911_ (.A0(_07254_),
    .A1(net2475),
    .S(_07231_),
    .X(_07255_));
 sky130_fd_sc_hd__clkbuf_1 _23912_ (.A(_07255_),
    .X(_02030_));
 sky130_fd_sc_hd__o211a_1 _23913_ (.A1(_12218_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07218_),
    .X(_07256_));
 sky130_fd_sc_hd__mux2_1 _23914_ (.A0(_07256_),
    .A1(net2411),
    .S(_07231_),
    .X(_07257_));
 sky130_fd_sc_hd__clkbuf_1 _23915_ (.A(_07257_),
    .X(_02031_));
 sky130_fd_sc_hd__o211a_1 _23916_ (.A1(_12226_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07221_),
    .X(_07258_));
 sky130_fd_sc_hd__mux2_1 _23917_ (.A0(_07258_),
    .A1(net2874),
    .S(_07231_),
    .X(_07259_));
 sky130_fd_sc_hd__clkbuf_1 _23918_ (.A(_07259_),
    .X(_02032_));
 sky130_fd_sc_hd__o211a_1 _23919_ (.A1(_12234_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07224_),
    .X(_07260_));
 sky130_fd_sc_hd__mux2_1 _23920_ (.A0(_07260_),
    .A1(net2834),
    .S(_07231_),
    .X(_07261_));
 sky130_fd_sc_hd__clkbuf_1 _23921_ (.A(_07261_),
    .X(_02033_));
 sky130_fd_sc_hd__o211a_1 _23922_ (.A1(_12242_),
    .A2(_07205_),
    .B1(_07247_),
    .C1(_07227_),
    .X(_07262_));
 sky130_fd_sc_hd__mux2_1 _23923_ (.A0(_07262_),
    .A1(net2337),
    .S(_07231_),
    .X(_07263_));
 sky130_fd_sc_hd__clkbuf_1 _23924_ (.A(_07263_),
    .X(_02034_));
 sky130_fd_sc_hd__nand2_1 _23925_ (.A(_07120_),
    .B(_04257_),
    .Y(_07264_));
 sky130_fd_sc_hd__a21bo_1 _23926_ (.A1(_07264_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_07265_));
 sky130_fd_sc_hd__clkbuf_8 _23927_ (.A(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__mux2_1 _23928_ (.A0(_06530_),
    .A1(net2396),
    .S(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__clkbuf_1 _23929_ (.A(_07267_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _23930_ (.A0(_06538_),
    .A1(net2584),
    .S(_07266_),
    .X(_07268_));
 sky130_fd_sc_hd__clkbuf_1 _23931_ (.A(_07268_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _23932_ (.A0(_06540_),
    .A1(net3390),
    .S(_07266_),
    .X(_07269_));
 sky130_fd_sc_hd__clkbuf_1 _23933_ (.A(_07269_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _23934_ (.A0(_06542_),
    .A1(net2631),
    .S(_07266_),
    .X(_07270_));
 sky130_fd_sc_hd__clkbuf_1 _23935_ (.A(_07270_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _23936_ (.A0(_06544_),
    .A1(net3055),
    .S(_07266_),
    .X(_07271_));
 sky130_fd_sc_hd__clkbuf_1 _23937_ (.A(_07271_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _23938_ (.A0(_06546_),
    .A1(net2941),
    .S(_07266_),
    .X(_07272_));
 sky130_fd_sc_hd__clkbuf_1 _23939_ (.A(_07272_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _23940_ (.A0(_06548_),
    .A1(net2819),
    .S(_07266_),
    .X(_07273_));
 sky130_fd_sc_hd__clkbuf_1 _23941_ (.A(_07273_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _23942_ (.A0(_06550_),
    .A1(net3527),
    .S(_07266_),
    .X(_07274_));
 sky130_fd_sc_hd__clkbuf_1 _23943_ (.A(_07274_),
    .X(_02042_));
 sky130_fd_sc_hd__buf_4 _23944_ (.A(_07264_),
    .X(_07275_));
 sky130_fd_sc_hd__buf_4 _23945_ (.A(_07264_),
    .X(_07276_));
 sky130_fd_sc_hd__nand2_1 _23946_ (.A(_07276_),
    .B(_12184_),
    .Y(_07277_));
 sky130_fd_sc_hd__o211a_1 _23947_ (.A1(_02850_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__mux2_1 _23948_ (.A0(_07278_),
    .A1(net2948),
    .S(_07266_),
    .X(_07279_));
 sky130_fd_sc_hd__clkbuf_1 _23949_ (.A(_07279_),
    .X(_02043_));
 sky130_fd_sc_hd__nand2_1 _23950_ (.A(_07276_),
    .B(_12197_),
    .Y(_07280_));
 sky130_fd_sc_hd__o211a_1 _23951_ (.A1(_02860_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__mux2_1 _23952_ (.A0(_07281_),
    .A1(net2296),
    .S(_07266_),
    .X(_07282_));
 sky130_fd_sc_hd__clkbuf_1 _23953_ (.A(_07282_),
    .X(_02044_));
 sky130_fd_sc_hd__nand2_1 _23954_ (.A(_07276_),
    .B(_12205_),
    .Y(_07283_));
 sky130_fd_sc_hd__o211a_1 _23955_ (.A1(_02867_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__mux2_1 _23956_ (.A0(_07284_),
    .A1(net2652),
    .S(_07266_),
    .X(_07285_));
 sky130_fd_sc_hd__clkbuf_1 _23957_ (.A(_07285_),
    .X(_02045_));
 sky130_fd_sc_hd__nand2_1 _23958_ (.A(_07276_),
    .B(_12213_),
    .Y(_07286_));
 sky130_fd_sc_hd__o211a_1 _23959_ (.A1(_02874_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__mux2_1 _23960_ (.A0(_07287_),
    .A1(net2746),
    .S(_07266_),
    .X(_07288_));
 sky130_fd_sc_hd__clkbuf_1 _23961_ (.A(_07288_),
    .X(_02046_));
 sky130_fd_sc_hd__nand2_1 _23962_ (.A(_07276_),
    .B(_12221_),
    .Y(_07289_));
 sky130_fd_sc_hd__o211a_1 _23963_ (.A1(_02881_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__mux2_1 _23964_ (.A0(_07290_),
    .A1(net3311),
    .S(_07266_),
    .X(_07291_));
 sky130_fd_sc_hd__clkbuf_1 _23965_ (.A(_07291_),
    .X(_02047_));
 sky130_fd_sc_hd__nand2_1 _23966_ (.A(_07276_),
    .B(_12229_),
    .Y(_07292_));
 sky130_fd_sc_hd__o211a_1 _23967_ (.A1(_02888_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__mux2_1 _23968_ (.A0(_07293_),
    .A1(net3408),
    .S(_07266_),
    .X(_07294_));
 sky130_fd_sc_hd__clkbuf_1 _23969_ (.A(_07294_),
    .X(_02048_));
 sky130_fd_sc_hd__nand2_1 _23970_ (.A(_07276_),
    .B(_12237_),
    .Y(_07295_));
 sky130_fd_sc_hd__o211a_1 _23971_ (.A1(_02895_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__mux2_1 _23972_ (.A0(_07296_),
    .A1(net3365),
    .S(_07266_),
    .X(_07297_));
 sky130_fd_sc_hd__clkbuf_1 _23973_ (.A(_07297_),
    .X(_02049_));
 sky130_fd_sc_hd__nand2_1 _23974_ (.A(_07276_),
    .B(_12245_),
    .Y(_07298_));
 sky130_fd_sc_hd__o211a_1 _23975_ (.A1(_02902_),
    .A2(_07275_),
    .B1(_07247_),
    .C1(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__mux2_1 _23976_ (.A0(_07299_),
    .A1(net2993),
    .S(_07266_),
    .X(_07300_));
 sky130_fd_sc_hd__clkbuf_1 _23977_ (.A(_07300_),
    .X(_02050_));
 sky130_fd_sc_hd__buf_4 _23978_ (.A(_06885_),
    .X(_07301_));
 sky130_fd_sc_hd__o211a_1 _23979_ (.A1(_02910_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07277_),
    .X(_07302_));
 sky130_fd_sc_hd__clkbuf_8 _23980_ (.A(_07265_),
    .X(_07303_));
 sky130_fd_sc_hd__mux2_1 _23981_ (.A0(_07302_),
    .A1(net3641),
    .S(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__clkbuf_1 _23982_ (.A(_07304_),
    .X(_02051_));
 sky130_fd_sc_hd__o211a_1 _23983_ (.A1(_02915_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07280_),
    .X(_07305_));
 sky130_fd_sc_hd__mux2_1 _23984_ (.A0(_07305_),
    .A1(net3473),
    .S(_07303_),
    .X(_07306_));
 sky130_fd_sc_hd__clkbuf_1 _23985_ (.A(_07306_),
    .X(_02052_));
 sky130_fd_sc_hd__o211a_1 _23986_ (.A1(_02920_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07283_),
    .X(_07307_));
 sky130_fd_sc_hd__mux2_1 _23987_ (.A0(_07307_),
    .A1(net2777),
    .S(_07303_),
    .X(_07308_));
 sky130_fd_sc_hd__clkbuf_1 _23988_ (.A(_07308_),
    .X(_02053_));
 sky130_fd_sc_hd__o211a_1 _23989_ (.A1(_02926_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07286_),
    .X(_07309_));
 sky130_fd_sc_hd__mux2_1 _23990_ (.A0(_07309_),
    .A1(net2841),
    .S(_07303_),
    .X(_07310_));
 sky130_fd_sc_hd__clkbuf_1 _23991_ (.A(_07310_),
    .X(_02054_));
 sky130_fd_sc_hd__o211a_1 _23992_ (.A1(_02931_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07289_),
    .X(_07311_));
 sky130_fd_sc_hd__mux2_1 _23993_ (.A0(_07311_),
    .A1(net2760),
    .S(_07303_),
    .X(_07312_));
 sky130_fd_sc_hd__clkbuf_1 _23994_ (.A(_07312_),
    .X(_02055_));
 sky130_fd_sc_hd__o211a_1 _23995_ (.A1(_02936_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07292_),
    .X(_07313_));
 sky130_fd_sc_hd__mux2_1 _23996_ (.A0(_07313_),
    .A1(net2508),
    .S(_07303_),
    .X(_07314_));
 sky130_fd_sc_hd__clkbuf_1 _23997_ (.A(_07314_),
    .X(_02056_));
 sky130_fd_sc_hd__o211a_1 _23998_ (.A1(_02941_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07295_),
    .X(_07315_));
 sky130_fd_sc_hd__mux2_1 _23999_ (.A0(_07315_),
    .A1(net3139),
    .S(_07303_),
    .X(_07316_));
 sky130_fd_sc_hd__clkbuf_1 _24000_ (.A(_07316_),
    .X(_02057_));
 sky130_fd_sc_hd__o211a_1 _24001_ (.A1(_02946_),
    .A2(_07275_),
    .B1(_07301_),
    .C1(_07298_),
    .X(_07317_));
 sky130_fd_sc_hd__mux2_1 _24002_ (.A0(_07317_),
    .A1(net3563),
    .S(_07303_),
    .X(_07318_));
 sky130_fd_sc_hd__clkbuf_1 _24003_ (.A(_07318_),
    .X(_02058_));
 sky130_fd_sc_hd__o211a_1 _24004_ (.A1(_12169_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07277_),
    .X(_07319_));
 sky130_fd_sc_hd__mux2_1 _24005_ (.A0(_07319_),
    .A1(net3097),
    .S(_07303_),
    .X(_07320_));
 sky130_fd_sc_hd__clkbuf_1 _24006_ (.A(_07320_),
    .X(_02059_));
 sky130_fd_sc_hd__o211a_1 _24007_ (.A1(_12194_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07280_),
    .X(_07321_));
 sky130_fd_sc_hd__mux2_1 _24008_ (.A0(_07321_),
    .A1(net3548),
    .S(_07303_),
    .X(_07322_));
 sky130_fd_sc_hd__clkbuf_1 _24009_ (.A(_07322_),
    .X(_02060_));
 sky130_fd_sc_hd__o211a_1 _24010_ (.A1(_12202_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07283_),
    .X(_07323_));
 sky130_fd_sc_hd__mux2_1 _24011_ (.A0(_07323_),
    .A1(net3720),
    .S(_07303_),
    .X(_07324_));
 sky130_fd_sc_hd__clkbuf_1 _24012_ (.A(_07324_),
    .X(_02061_));
 sky130_fd_sc_hd__o211a_1 _24013_ (.A1(_12210_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07286_),
    .X(_07325_));
 sky130_fd_sc_hd__mux2_1 _24014_ (.A0(_07325_),
    .A1(net3708),
    .S(_07303_),
    .X(_07326_));
 sky130_fd_sc_hd__clkbuf_1 _24015_ (.A(_07326_),
    .X(_02062_));
 sky130_fd_sc_hd__o211a_1 _24016_ (.A1(_12218_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07289_),
    .X(_07327_));
 sky130_fd_sc_hd__mux2_1 _24017_ (.A0(_07327_),
    .A1(net3787),
    .S(_07303_),
    .X(_07328_));
 sky130_fd_sc_hd__clkbuf_1 _24018_ (.A(_07328_),
    .X(_02063_));
 sky130_fd_sc_hd__o211a_1 _24019_ (.A1(_12226_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07292_),
    .X(_07329_));
 sky130_fd_sc_hd__mux2_1 _24020_ (.A0(_07329_),
    .A1(net3795),
    .S(_07303_),
    .X(_07330_));
 sky130_fd_sc_hd__clkbuf_1 _24021_ (.A(_07330_),
    .X(_02064_));
 sky130_fd_sc_hd__o211a_1 _24022_ (.A1(_12234_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07295_),
    .X(_07331_));
 sky130_fd_sc_hd__mux2_1 _24023_ (.A0(_07331_),
    .A1(net3751),
    .S(_07303_),
    .X(_07332_));
 sky130_fd_sc_hd__clkbuf_1 _24024_ (.A(_07332_),
    .X(_02065_));
 sky130_fd_sc_hd__o211a_1 _24025_ (.A1(_12242_),
    .A2(_07276_),
    .B1(_07301_),
    .C1(_07298_),
    .X(_07333_));
 sky130_fd_sc_hd__mux2_1 _24026_ (.A0(_07333_),
    .A1(net3653),
    .S(_07303_),
    .X(_07334_));
 sky130_fd_sc_hd__clkbuf_1 _24027_ (.A(_07334_),
    .X(_02066_));
 sky130_fd_sc_hd__nand2_1 _24028_ (.A(_07120_),
    .B(_04333_),
    .Y(_07335_));
 sky130_fd_sc_hd__inv_2 _24029_ (.A(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__o21ai_4 _24030_ (.A1(_06755_),
    .A2(_07336_),
    .B1(_06020_),
    .Y(_07337_));
 sky130_fd_sc_hd__mux2_1 _24031_ (.A0(_06530_),
    .A1(net2773),
    .S(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__clkbuf_1 _24032_ (.A(_07338_),
    .X(_02067_));
 sky130_fd_sc_hd__mux2_1 _24033_ (.A0(_06538_),
    .A1(net2355),
    .S(_07337_),
    .X(_07339_));
 sky130_fd_sc_hd__clkbuf_1 _24034_ (.A(_07339_),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _24035_ (.A0(_06540_),
    .A1(net3177),
    .S(_07337_),
    .X(_07340_));
 sky130_fd_sc_hd__clkbuf_1 _24036_ (.A(_07340_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _24037_ (.A0(_06542_),
    .A1(net3103),
    .S(_07337_),
    .X(_07341_));
 sky130_fd_sc_hd__clkbuf_1 _24038_ (.A(_07341_),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _24039_ (.A0(_06544_),
    .A1(net3363),
    .S(_07337_),
    .X(_07342_));
 sky130_fd_sc_hd__clkbuf_1 _24040_ (.A(_07342_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _24041_ (.A0(_06546_),
    .A1(net2156),
    .S(_07337_),
    .X(_07343_));
 sky130_fd_sc_hd__clkbuf_1 _24042_ (.A(_07343_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _24043_ (.A0(_06548_),
    .A1(net2636),
    .S(_07337_),
    .X(_07344_));
 sky130_fd_sc_hd__clkbuf_1 _24044_ (.A(_07344_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _24045_ (.A0(_06550_),
    .A1(net3134),
    .S(_07337_),
    .X(_07345_));
 sky130_fd_sc_hd__clkbuf_1 _24046_ (.A(_07345_),
    .X(_02074_));
 sky130_fd_sc_hd__buf_4 _24047_ (.A(_07337_),
    .X(_07346_));
 sky130_fd_sc_hd__buf_4 _24048_ (.A(_07336_),
    .X(_07347_));
 sky130_fd_sc_hd__buf_4 _24049_ (.A(_07336_),
    .X(_07348_));
 sky130_fd_sc_hd__nor2_1 _24050_ (.A(_05583_),
    .B(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__a211o_1 _24051_ (.A1(_05484_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__buf_4 _24052_ (.A(_07337_),
    .X(_07351_));
 sky130_fd_sc_hd__nand2_1 _24053_ (.A(_07351_),
    .B(net1010),
    .Y(_07352_));
 sky130_fd_sc_hd__o21ai_1 _24054_ (.A1(_07346_),
    .A2(_07350_),
    .B1(net1011),
    .Y(_02075_));
 sky130_fd_sc_hd__nor2_1 _24055_ (.A(_05589_),
    .B(_07348_),
    .Y(_07353_));
 sky130_fd_sc_hd__a211o_1 _24056_ (.A1(_05491_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__nand2_1 _24057_ (.A(_07351_),
    .B(net852),
    .Y(_07355_));
 sky130_fd_sc_hd__o21ai_1 _24058_ (.A1(_07346_),
    .A2(_07354_),
    .B1(net853),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _24059_ (.A(_05593_),
    .B(_07348_),
    .Y(_07356_));
 sky130_fd_sc_hd__a211o_1 _24060_ (.A1(_05495_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__nand2_1 _24061_ (.A(_07351_),
    .B(net1004),
    .Y(_07358_));
 sky130_fd_sc_hd__o21ai_1 _24062_ (.A1(_07346_),
    .A2(_07357_),
    .B1(net1005),
    .Y(_02077_));
 sky130_fd_sc_hd__nor2_1 _24063_ (.A(_05597_),
    .B(_07348_),
    .Y(_07359_));
 sky130_fd_sc_hd__a211o_1 _24064_ (.A1(_05500_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07359_),
    .X(_07360_));
 sky130_fd_sc_hd__nand2_1 _24065_ (.A(_07351_),
    .B(net1130),
    .Y(_07361_));
 sky130_fd_sc_hd__o21ai_1 _24066_ (.A1(_07346_),
    .A2(_07360_),
    .B1(net1131),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _24067_ (.A(_05601_),
    .B(_07348_),
    .Y(_07362_));
 sky130_fd_sc_hd__a211o_1 _24068_ (.A1(_05504_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__nand2_1 _24069_ (.A(_07351_),
    .B(net1871),
    .Y(_07364_));
 sky130_fd_sc_hd__o21ai_1 _24070_ (.A1(_07346_),
    .A2(_07363_),
    .B1(net1872),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _24071_ (.A(_05605_),
    .B(_07348_),
    .Y(_07365_));
 sky130_fd_sc_hd__a211o_1 _24072_ (.A1(_05508_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07365_),
    .X(_07366_));
 sky130_fd_sc_hd__nand2_1 _24073_ (.A(_07351_),
    .B(net860),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_1 _24074_ (.A1(_07346_),
    .A2(_07366_),
    .B1(net861),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _24075_ (.A(_05609_),
    .B(_07348_),
    .Y(_07368_));
 sky130_fd_sc_hd__a211o_1 _24076_ (.A1(_05512_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07368_),
    .X(_07369_));
 sky130_fd_sc_hd__nand2_1 _24077_ (.A(_07351_),
    .B(net1370),
    .Y(_07370_));
 sky130_fd_sc_hd__o21ai_1 _24078_ (.A1(_07346_),
    .A2(_07369_),
    .B1(net1371),
    .Y(_02081_));
 sky130_fd_sc_hd__nor2_1 _24079_ (.A(_05613_),
    .B(_07348_),
    .Y(_07371_));
 sky130_fd_sc_hd__a211o_1 _24080_ (.A1(_05516_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(_07351_),
    .B(net1734),
    .Y(_07373_));
 sky130_fd_sc_hd__o21ai_1 _24082_ (.A1(_07346_),
    .A2(_07372_),
    .B1(net1735),
    .Y(_02082_));
 sky130_fd_sc_hd__buf_4 _24083_ (.A(_07337_),
    .X(_07374_));
 sky130_fd_sc_hd__a211o_1 _24084_ (.A1(_05521_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07349_),
    .X(_07375_));
 sky130_fd_sc_hd__nand2_1 _24085_ (.A(_07351_),
    .B(net1544),
    .Y(_07376_));
 sky130_fd_sc_hd__o21ai_1 _24086_ (.A1(_07374_),
    .A2(_07375_),
    .B1(net1545),
    .Y(_02083_));
 sky130_fd_sc_hd__a211o_1 _24087_ (.A1(_05524_),
    .A2(_07347_),
    .B1(_07107_),
    .C1(_07353_),
    .X(_07377_));
 sky130_fd_sc_hd__nand2_1 _24088_ (.A(_07351_),
    .B(net1394),
    .Y(_07378_));
 sky130_fd_sc_hd__o21ai_1 _24089_ (.A1(_07374_),
    .A2(_07377_),
    .B1(net1395),
    .Y(_02084_));
 sky130_fd_sc_hd__buf_4 _24090_ (.A(_05892_),
    .X(_07379_));
 sky130_fd_sc_hd__a211o_1 _24091_ (.A1(_05527_),
    .A2(_07347_),
    .B1(_07379_),
    .C1(_07356_),
    .X(_07380_));
 sky130_fd_sc_hd__nand2_1 _24092_ (.A(_07351_),
    .B(net1708),
    .Y(_07381_));
 sky130_fd_sc_hd__o21ai_1 _24093_ (.A1(_07374_),
    .A2(_07380_),
    .B1(net1709),
    .Y(_02085_));
 sky130_fd_sc_hd__a211o_1 _24094_ (.A1(_05530_),
    .A2(_07347_),
    .B1(_07379_),
    .C1(_07359_),
    .X(_07382_));
 sky130_fd_sc_hd__nand2_1 _24095_ (.A(_07351_),
    .B(net1684),
    .Y(_07383_));
 sky130_fd_sc_hd__o21ai_1 _24096_ (.A1(_07374_),
    .A2(_07382_),
    .B1(net1685),
    .Y(_02086_));
 sky130_fd_sc_hd__a211o_1 _24097_ (.A1(_05533_),
    .A2(_07347_),
    .B1(_07379_),
    .C1(_07362_),
    .X(_07384_));
 sky130_fd_sc_hd__nand2_1 _24098_ (.A(_07351_),
    .B(net1076),
    .Y(_07385_));
 sky130_fd_sc_hd__o21ai_1 _24099_ (.A1(_07374_),
    .A2(_07384_),
    .B1(net1077),
    .Y(_02087_));
 sky130_fd_sc_hd__a211o_1 _24100_ (.A1(_05536_),
    .A2(_07347_),
    .B1(_07379_),
    .C1(_07365_),
    .X(_07386_));
 sky130_fd_sc_hd__nand2_1 _24101_ (.A(_07351_),
    .B(net1418),
    .Y(_07387_));
 sky130_fd_sc_hd__o21ai_1 _24102_ (.A1(_07374_),
    .A2(_07386_),
    .B1(net1419),
    .Y(_02088_));
 sky130_fd_sc_hd__a211o_1 _24103_ (.A1(_05539_),
    .A2(_07347_),
    .B1(_07379_),
    .C1(_07368_),
    .X(_07388_));
 sky130_fd_sc_hd__nand2_1 _24104_ (.A(_07351_),
    .B(net740),
    .Y(_07389_));
 sky130_fd_sc_hd__o21ai_1 _24105_ (.A1(_07374_),
    .A2(_07388_),
    .B1(net741),
    .Y(_02089_));
 sky130_fd_sc_hd__a211o_1 _24106_ (.A1(_05542_),
    .A2(_07347_),
    .B1(_07379_),
    .C1(_07371_),
    .X(_07390_));
 sky130_fd_sc_hd__nand2_1 _24107_ (.A(_07351_),
    .B(net1818),
    .Y(_07391_));
 sky130_fd_sc_hd__o21ai_1 _24108_ (.A1(_07374_),
    .A2(_07390_),
    .B1(net1819),
    .Y(_02090_));
 sky130_fd_sc_hd__a211o_1 _24109_ (.A1(_05545_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07349_),
    .X(_07392_));
 sky130_fd_sc_hd__nand2_1 _24110_ (.A(_07346_),
    .B(net1722),
    .Y(_07393_));
 sky130_fd_sc_hd__o21ai_1 _24111_ (.A1(_07374_),
    .A2(_07392_),
    .B1(net1723),
    .Y(_02091_));
 sky130_fd_sc_hd__a211o_1 _24112_ (.A1(_05548_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07353_),
    .X(_07394_));
 sky130_fd_sc_hd__nand2_1 _24113_ (.A(_07346_),
    .B(net1816),
    .Y(_07395_));
 sky130_fd_sc_hd__o21ai_1 _24114_ (.A1(_07374_),
    .A2(_07394_),
    .B1(net1817),
    .Y(_02092_));
 sky130_fd_sc_hd__a211o_1 _24115_ (.A1(_05551_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07356_),
    .X(_07396_));
 sky130_fd_sc_hd__nand2_1 _24116_ (.A(_07346_),
    .B(net1350),
    .Y(_07397_));
 sky130_fd_sc_hd__o21ai_1 _24117_ (.A1(_07374_),
    .A2(_07396_),
    .B1(net1351),
    .Y(_02093_));
 sky130_fd_sc_hd__a211o_1 _24118_ (.A1(_05555_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07359_),
    .X(_07398_));
 sky130_fd_sc_hd__nand2_1 _24119_ (.A(_07346_),
    .B(net1538),
    .Y(_07399_));
 sky130_fd_sc_hd__o21ai_1 _24120_ (.A1(_07374_),
    .A2(_07398_),
    .B1(net1539),
    .Y(_02094_));
 sky130_fd_sc_hd__a211o_1 _24121_ (.A1(_05558_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07362_),
    .X(_07400_));
 sky130_fd_sc_hd__nand2_1 _24122_ (.A(_07346_),
    .B(net1546),
    .Y(_07401_));
 sky130_fd_sc_hd__o21ai_1 _24123_ (.A1(_07374_),
    .A2(_07400_),
    .B1(net1547),
    .Y(_02095_));
 sky130_fd_sc_hd__a211o_1 _24124_ (.A1(_05561_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07365_),
    .X(_07402_));
 sky130_fd_sc_hd__nand2_1 _24125_ (.A(_07346_),
    .B(net1124),
    .Y(_07403_));
 sky130_fd_sc_hd__o21ai_1 _24126_ (.A1(_07374_),
    .A2(_07402_),
    .B1(net1125),
    .Y(_02096_));
 sky130_fd_sc_hd__a211o_1 _24127_ (.A1(_05564_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07368_),
    .X(_07404_));
 sky130_fd_sc_hd__nand2_1 _24128_ (.A(_07346_),
    .B(net1800),
    .Y(_07405_));
 sky130_fd_sc_hd__o21ai_1 _24129_ (.A1(_07374_),
    .A2(_07404_),
    .B1(net1801),
    .Y(_02097_));
 sky130_fd_sc_hd__a211o_1 _24130_ (.A1(_05567_),
    .A2(_07348_),
    .B1(_07379_),
    .C1(_07371_),
    .X(_07406_));
 sky130_fd_sc_hd__nand2_1 _24131_ (.A(_07346_),
    .B(net1934),
    .Y(_07407_));
 sky130_fd_sc_hd__o21ai_1 _24132_ (.A1(_07374_),
    .A2(_07406_),
    .B1(_07407_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand2_1 _24133_ (.A(_04104_),
    .B(_12311_),
    .Y(_07408_));
 sky130_fd_sc_hd__inv_2 _24134_ (.A(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__o21ai_4 _24135_ (.A1(_06755_),
    .A2(_07409_),
    .B1(_06020_),
    .Y(_07410_));
 sky130_fd_sc_hd__mux2_1 _24136_ (.A0(_06530_),
    .A1(net2375),
    .S(_07410_),
    .X(_07411_));
 sky130_fd_sc_hd__clkbuf_1 _24137_ (.A(_07411_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _24138_ (.A0(_06538_),
    .A1(net3138),
    .S(_07410_),
    .X(_07412_));
 sky130_fd_sc_hd__clkbuf_1 _24139_ (.A(_07412_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _24140_ (.A0(_06540_),
    .A1(net2724),
    .S(_07410_),
    .X(_07413_));
 sky130_fd_sc_hd__clkbuf_1 _24141_ (.A(_07413_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _24142_ (.A0(_06542_),
    .A1(net2447),
    .S(_07410_),
    .X(_07414_));
 sky130_fd_sc_hd__clkbuf_1 _24143_ (.A(_07414_),
    .X(_02102_));
 sky130_fd_sc_hd__mux2_1 _24144_ (.A0(_06544_),
    .A1(net2123),
    .S(_07410_),
    .X(_07415_));
 sky130_fd_sc_hd__clkbuf_1 _24145_ (.A(_07415_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _24146_ (.A0(_06546_),
    .A1(net2048),
    .S(_07410_),
    .X(_07416_));
 sky130_fd_sc_hd__clkbuf_1 _24147_ (.A(_07416_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _24148_ (.A0(_06548_),
    .A1(net2114),
    .S(_07410_),
    .X(_07417_));
 sky130_fd_sc_hd__clkbuf_1 _24149_ (.A(_07417_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _24150_ (.A0(_06550_),
    .A1(net2367),
    .S(_07410_),
    .X(_07418_));
 sky130_fd_sc_hd__clkbuf_1 _24151_ (.A(_07418_),
    .X(_02106_));
 sky130_fd_sc_hd__buf_4 _24152_ (.A(_07410_),
    .X(_07419_));
 sky130_fd_sc_hd__buf_4 _24153_ (.A(_07409_),
    .X(_07420_));
 sky130_fd_sc_hd__buf_4 _24154_ (.A(_07409_),
    .X(_07421_));
 sky130_fd_sc_hd__nor2_1 _24155_ (.A(_05583_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__a211o_1 _24156_ (.A1(_05484_),
    .A2(_07420_),
    .B1(_07379_),
    .C1(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__buf_4 _24157_ (.A(_07410_),
    .X(_07424_));
 sky130_fd_sc_hd__nand2_1 _24158_ (.A(_07424_),
    .B(net1172),
    .Y(_07425_));
 sky130_fd_sc_hd__o21ai_1 _24159_ (.A1(_07419_),
    .A2(_07423_),
    .B1(net1173),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_1 _24160_ (.A(_05589_),
    .B(_07421_),
    .Y(_07426_));
 sky130_fd_sc_hd__a211o_1 _24161_ (.A1(_05491_),
    .A2(_07420_),
    .B1(_07379_),
    .C1(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__nand2_1 _24162_ (.A(_07424_),
    .B(net492),
    .Y(_07428_));
 sky130_fd_sc_hd__o21ai_1 _24163_ (.A1(_07419_),
    .A2(_07427_),
    .B1(net493),
    .Y(_02108_));
 sky130_fd_sc_hd__buf_4 _24164_ (.A(_05892_),
    .X(_07429_));
 sky130_fd_sc_hd__nor2_1 _24165_ (.A(_05593_),
    .B(_07421_),
    .Y(_07430_));
 sky130_fd_sc_hd__a211o_1 _24166_ (.A1(_05495_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__nand2_1 _24167_ (.A(_07424_),
    .B(net1932),
    .Y(_07432_));
 sky130_fd_sc_hd__o21ai_1 _24168_ (.A1(_07419_),
    .A2(_07431_),
    .B1(net1933),
    .Y(_02109_));
 sky130_fd_sc_hd__nor2_1 _24169_ (.A(_05597_),
    .B(_07421_),
    .Y(_07433_));
 sky130_fd_sc_hd__a211o_1 _24170_ (.A1(_05500_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__nand2_1 _24171_ (.A(_07424_),
    .B(net1634),
    .Y(_07435_));
 sky130_fd_sc_hd__o21ai_1 _24172_ (.A1(_07419_),
    .A2(_07434_),
    .B1(net1635),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_1 _24173_ (.A(_05601_),
    .B(_07421_),
    .Y(_07436_));
 sky130_fd_sc_hd__a211o_1 _24174_ (.A1(_05504_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__nand2_1 _24175_ (.A(_07424_),
    .B(net478),
    .Y(_07438_));
 sky130_fd_sc_hd__o21ai_1 _24176_ (.A1(_07419_),
    .A2(_07437_),
    .B1(net479),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _24177_ (.A(_05605_),
    .B(_07421_),
    .Y(_07439_));
 sky130_fd_sc_hd__a211o_1 _24178_ (.A1(_05508_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__nand2_1 _24179_ (.A(_07424_),
    .B(net1846),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_1 _24180_ (.A1(_07419_),
    .A2(_07440_),
    .B1(net1847),
    .Y(_02112_));
 sky130_fd_sc_hd__nor2_1 _24181_ (.A(_05609_),
    .B(_07421_),
    .Y(_07442_));
 sky130_fd_sc_hd__a211o_1 _24182_ (.A1(_05512_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__nand2_1 _24183_ (.A(_07424_),
    .B(net1961),
    .Y(_07444_));
 sky130_fd_sc_hd__o21ai_1 _24184_ (.A1(_07419_),
    .A2(_07443_),
    .B1(_07444_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _24185_ (.A(_05613_),
    .B(_07421_),
    .Y(_07445_));
 sky130_fd_sc_hd__a211o_1 _24186_ (.A1(_05516_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__nand2_1 _24187_ (.A(_07424_),
    .B(net520),
    .Y(_07447_));
 sky130_fd_sc_hd__o21ai_1 _24188_ (.A1(_07419_),
    .A2(_07446_),
    .B1(net521),
    .Y(_02114_));
 sky130_fd_sc_hd__buf_4 _24189_ (.A(_07410_),
    .X(_07448_));
 sky130_fd_sc_hd__a211o_1 _24190_ (.A1(_05521_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07422_),
    .X(_07449_));
 sky130_fd_sc_hd__nand2_1 _24191_ (.A(_07424_),
    .B(net1834),
    .Y(_07450_));
 sky130_fd_sc_hd__o21ai_1 _24192_ (.A1(_07448_),
    .A2(_07449_),
    .B1(net1835),
    .Y(_02115_));
 sky130_fd_sc_hd__a211o_1 _24193_ (.A1(_05524_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07426_),
    .X(_07451_));
 sky130_fd_sc_hd__nand2_1 _24194_ (.A(_07424_),
    .B(net1973),
    .Y(_07452_));
 sky130_fd_sc_hd__o21ai_1 _24195_ (.A1(_07448_),
    .A2(_07451_),
    .B1(_07452_),
    .Y(_02116_));
 sky130_fd_sc_hd__a211o_1 _24196_ (.A1(_05527_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07430_),
    .X(_07453_));
 sky130_fd_sc_hd__nand2_1 _24197_ (.A(_07424_),
    .B(net1969),
    .Y(_07454_));
 sky130_fd_sc_hd__o21ai_1 _24198_ (.A1(_07448_),
    .A2(_07453_),
    .B1(_07454_),
    .Y(_02117_));
 sky130_fd_sc_hd__a211o_1 _24199_ (.A1(_05530_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07433_),
    .X(_07455_));
 sky130_fd_sc_hd__nand2_1 _24200_ (.A(_07424_),
    .B(net1276),
    .Y(_07456_));
 sky130_fd_sc_hd__o21ai_1 _24201_ (.A1(_07448_),
    .A2(_07455_),
    .B1(net1277),
    .Y(_02118_));
 sky130_fd_sc_hd__a211o_1 _24202_ (.A1(_05533_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07436_),
    .X(_07457_));
 sky130_fd_sc_hd__nand2_1 _24203_ (.A(_07424_),
    .B(net594),
    .Y(_07458_));
 sky130_fd_sc_hd__o21ai_1 _24204_ (.A1(_07448_),
    .A2(_07457_),
    .B1(net595),
    .Y(_02119_));
 sky130_fd_sc_hd__a211o_1 _24205_ (.A1(_05536_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07439_),
    .X(_07459_));
 sky130_fd_sc_hd__nand2_1 _24206_ (.A(_07424_),
    .B(net1188),
    .Y(_07460_));
 sky130_fd_sc_hd__o21ai_1 _24207_ (.A1(_07448_),
    .A2(_07459_),
    .B1(net1189),
    .Y(_02120_));
 sky130_fd_sc_hd__a211o_1 _24208_ (.A1(_05539_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07442_),
    .X(_07461_));
 sky130_fd_sc_hd__nand2_1 _24209_ (.A(_07424_),
    .B(net1980),
    .Y(_07462_));
 sky130_fd_sc_hd__o21ai_1 _24210_ (.A1(_07448_),
    .A2(_07461_),
    .B1(_07462_),
    .Y(_02121_));
 sky130_fd_sc_hd__a211o_1 _24211_ (.A1(_05542_),
    .A2(_07420_),
    .B1(_07429_),
    .C1(_07445_),
    .X(_07463_));
 sky130_fd_sc_hd__nand2_1 _24212_ (.A(_07424_),
    .B(net1568),
    .Y(_07464_));
 sky130_fd_sc_hd__o21ai_1 _24213_ (.A1(_07448_),
    .A2(_07463_),
    .B1(net1569),
    .Y(_02122_));
 sky130_fd_sc_hd__a211o_1 _24214_ (.A1(_05545_),
    .A2(_07421_),
    .B1(_07429_),
    .C1(_07422_),
    .X(_07465_));
 sky130_fd_sc_hd__nand2_1 _24215_ (.A(_07419_),
    .B(net1869),
    .Y(_07466_));
 sky130_fd_sc_hd__o21ai_1 _24216_ (.A1(_07448_),
    .A2(_07465_),
    .B1(net1870),
    .Y(_02123_));
 sky130_fd_sc_hd__a211o_1 _24217_ (.A1(_05548_),
    .A2(_07421_),
    .B1(_07429_),
    .C1(_07426_),
    .X(_07467_));
 sky130_fd_sc_hd__nand2_1 _24218_ (.A(_07419_),
    .B(net1891),
    .Y(_07468_));
 sky130_fd_sc_hd__o21ai_1 _24219_ (.A1(_07448_),
    .A2(_07467_),
    .B1(net1892),
    .Y(_02124_));
 sky130_fd_sc_hd__buf_4 _24220_ (.A(_05892_),
    .X(_07469_));
 sky130_fd_sc_hd__a211o_1 _24221_ (.A1(_05551_),
    .A2(_07421_),
    .B1(_07469_),
    .C1(_07430_),
    .X(_07470_));
 sky130_fd_sc_hd__nand2_1 _24222_ (.A(_07419_),
    .B(net1754),
    .Y(_07471_));
 sky130_fd_sc_hd__o21ai_1 _24223_ (.A1(_07448_),
    .A2(_07470_),
    .B1(net1755),
    .Y(_02125_));
 sky130_fd_sc_hd__a211o_1 _24224_ (.A1(_05555_),
    .A2(_07421_),
    .B1(_07469_),
    .C1(_07433_),
    .X(_07472_));
 sky130_fd_sc_hd__nand2_1 _24225_ (.A(_07419_),
    .B(net442),
    .Y(_07473_));
 sky130_fd_sc_hd__o21ai_1 _24226_ (.A1(_07448_),
    .A2(_07472_),
    .B1(net443),
    .Y(_02126_));
 sky130_fd_sc_hd__a211o_1 _24227_ (.A1(_05558_),
    .A2(_07421_),
    .B1(_07469_),
    .C1(_07436_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_1 _24228_ (.A(_07419_),
    .B(net428),
    .Y(_07475_));
 sky130_fd_sc_hd__o21ai_1 _24229_ (.A1(_07448_),
    .A2(_07474_),
    .B1(net429),
    .Y(_02127_));
 sky130_fd_sc_hd__a211o_1 _24230_ (.A1(_05561_),
    .A2(_07421_),
    .B1(_07469_),
    .C1(_07439_),
    .X(_07476_));
 sky130_fd_sc_hd__nand2_1 _24231_ (.A(_07419_),
    .B(net420),
    .Y(_07477_));
 sky130_fd_sc_hd__o21ai_1 _24232_ (.A1(_07448_),
    .A2(_07476_),
    .B1(net421),
    .Y(_02128_));
 sky130_fd_sc_hd__a211o_1 _24233_ (.A1(_05564_),
    .A2(_07421_),
    .B1(_07469_),
    .C1(_07442_),
    .X(_07478_));
 sky130_fd_sc_hd__nand2_1 _24234_ (.A(_07419_),
    .B(net758),
    .Y(_07479_));
 sky130_fd_sc_hd__o21ai_1 _24235_ (.A1(_07448_),
    .A2(_07478_),
    .B1(net759),
    .Y(_02129_));
 sky130_fd_sc_hd__a211o_1 _24236_ (.A1(_05567_),
    .A2(_07421_),
    .B1(_07469_),
    .C1(_07445_),
    .X(_07480_));
 sky130_fd_sc_hd__nand2_1 _24237_ (.A(_07419_),
    .B(net588),
    .Y(_07481_));
 sky130_fd_sc_hd__o21ai_1 _24238_ (.A1(_07448_),
    .A2(_07480_),
    .B1(net589),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _24239_ (.A(_04183_),
    .B(_12311_),
    .Y(_07482_));
 sky130_fd_sc_hd__inv_2 _24240_ (.A(_07482_),
    .Y(_07483_));
 sky130_fd_sc_hd__o21ai_4 _24241_ (.A1(_06755_),
    .A2(_07483_),
    .B1(_06020_),
    .Y(_07484_));
 sky130_fd_sc_hd__mux2_1 _24242_ (.A0(_06530_),
    .A1(net2212),
    .S(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__clkbuf_1 _24243_ (.A(_07485_),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _24244_ (.A0(_06538_),
    .A1(net2153),
    .S(_07484_),
    .X(_07486_));
 sky130_fd_sc_hd__clkbuf_1 _24245_ (.A(_07486_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _24246_ (.A0(_06540_),
    .A1(net2109),
    .S(_07484_),
    .X(_07487_));
 sky130_fd_sc_hd__clkbuf_1 _24247_ (.A(_07487_),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _24248_ (.A0(_06542_),
    .A1(net2055),
    .S(_07484_),
    .X(_07488_));
 sky130_fd_sc_hd__clkbuf_1 _24249_ (.A(_07488_),
    .X(_02134_));
 sky130_fd_sc_hd__mux2_1 _24250_ (.A0(_06544_),
    .A1(net2119),
    .S(_07484_),
    .X(_07489_));
 sky130_fd_sc_hd__clkbuf_1 _24251_ (.A(_07489_),
    .X(_02135_));
 sky130_fd_sc_hd__mux2_1 _24252_ (.A0(_06546_),
    .A1(net2083),
    .S(_07484_),
    .X(_07490_));
 sky130_fd_sc_hd__clkbuf_1 _24253_ (.A(_07490_),
    .X(_02136_));
 sky130_fd_sc_hd__mux2_1 _24254_ (.A0(_06548_),
    .A1(net2041),
    .S(_07484_),
    .X(_07491_));
 sky130_fd_sc_hd__clkbuf_1 _24255_ (.A(_07491_),
    .X(_02137_));
 sky130_fd_sc_hd__mux2_1 _24256_ (.A0(_06550_),
    .A1(net2032),
    .S(_07484_),
    .X(_07492_));
 sky130_fd_sc_hd__clkbuf_1 _24257_ (.A(_07492_),
    .X(_02138_));
 sky130_fd_sc_hd__buf_4 _24258_ (.A(_07484_),
    .X(_07493_));
 sky130_fd_sc_hd__buf_4 _24259_ (.A(_07483_),
    .X(_07494_));
 sky130_fd_sc_hd__buf_4 _24260_ (.A(_07483_),
    .X(_07495_));
 sky130_fd_sc_hd__nor2_1 _24261_ (.A(_05583_),
    .B(_07495_),
    .Y(_07496_));
 sky130_fd_sc_hd__a211o_1 _24262_ (.A1(_05484_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__buf_4 _24263_ (.A(_07484_),
    .X(_07498_));
 sky130_fd_sc_hd__nand2_1 _24264_ (.A(_07498_),
    .B(net582),
    .Y(_07499_));
 sky130_fd_sc_hd__o21ai_1 _24265_ (.A1(_07493_),
    .A2(_07497_),
    .B1(net583),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_1 _24266_ (.A(_05589_),
    .B(_07495_),
    .Y(_07500_));
 sky130_fd_sc_hd__a211o_1 _24267_ (.A1(_05491_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__nand2_1 _24268_ (.A(_07498_),
    .B(net1558),
    .Y(_07502_));
 sky130_fd_sc_hd__o21ai_1 _24269_ (.A1(_07493_),
    .A2(_07501_),
    .B1(net1559),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _24270_ (.A(_05593_),
    .B(_07495_),
    .Y(_07503_));
 sky130_fd_sc_hd__a211o_1 _24271_ (.A1(_05495_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__nand2_1 _24272_ (.A(_07498_),
    .B(net1780),
    .Y(_07505_));
 sky130_fd_sc_hd__o21ai_1 _24273_ (.A1(_07493_),
    .A2(_07504_),
    .B1(net1781),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_1 _24274_ (.A(_05597_),
    .B(_07495_),
    .Y(_07506_));
 sky130_fd_sc_hd__a211o_1 _24275_ (.A1(_05500_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07506_),
    .X(_07507_));
 sky130_fd_sc_hd__nand2_1 _24276_ (.A(_07498_),
    .B(net476),
    .Y(_07508_));
 sky130_fd_sc_hd__o21ai_1 _24277_ (.A1(_07493_),
    .A2(_07507_),
    .B1(net477),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _24278_ (.A(_05601_),
    .B(_07495_),
    .Y(_07509_));
 sky130_fd_sc_hd__a211o_1 _24279_ (.A1(_05504_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__nand2_1 _24280_ (.A(_07498_),
    .B(net496),
    .Y(_07511_));
 sky130_fd_sc_hd__o21ai_1 _24281_ (.A1(_07493_),
    .A2(_07510_),
    .B1(net497),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _24282_ (.A(_05605_),
    .B(_07495_),
    .Y(_07512_));
 sky130_fd_sc_hd__a211o_1 _24283_ (.A1(_05508_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__nand2_1 _24284_ (.A(_07498_),
    .B(net1232),
    .Y(_07514_));
 sky130_fd_sc_hd__o21ai_1 _24285_ (.A1(_07493_),
    .A2(_07513_),
    .B1(net1233),
    .Y(_02144_));
 sky130_fd_sc_hd__nor2_1 _24286_ (.A(_05609_),
    .B(_07495_),
    .Y(_07515_));
 sky130_fd_sc_hd__a211o_1 _24287_ (.A1(_05512_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__nand2_1 _24288_ (.A(_07498_),
    .B(net628),
    .Y(_07517_));
 sky130_fd_sc_hd__o21ai_1 _24289_ (.A1(_07493_),
    .A2(_07516_),
    .B1(net629),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _24290_ (.A(_05613_),
    .B(_07495_),
    .Y(_07518_));
 sky130_fd_sc_hd__a211o_1 _24291_ (.A1(_05516_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07518_),
    .X(_07519_));
 sky130_fd_sc_hd__nand2_1 _24292_ (.A(_07498_),
    .B(net546),
    .Y(_07520_));
 sky130_fd_sc_hd__o21ai_1 _24293_ (.A1(_07493_),
    .A2(_07519_),
    .B1(net547),
    .Y(_02146_));
 sky130_fd_sc_hd__buf_4 _24294_ (.A(_07484_),
    .X(_07521_));
 sky130_fd_sc_hd__a211o_1 _24295_ (.A1(_05521_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07496_),
    .X(_07522_));
 sky130_fd_sc_hd__nand2_1 _24296_ (.A(_07498_),
    .B(net618),
    .Y(_07523_));
 sky130_fd_sc_hd__o21ai_1 _24297_ (.A1(_07521_),
    .A2(_07522_),
    .B1(net619),
    .Y(_02147_));
 sky130_fd_sc_hd__a211o_1 _24298_ (.A1(_05524_),
    .A2(_07494_),
    .B1(_07469_),
    .C1(_07500_),
    .X(_07524_));
 sky130_fd_sc_hd__nand2_1 _24299_ (.A(_07498_),
    .B(net458),
    .Y(_07525_));
 sky130_fd_sc_hd__o21ai_1 _24300_ (.A1(_07521_),
    .A2(_07524_),
    .B1(net459),
    .Y(_02148_));
 sky130_fd_sc_hd__buf_4 _24301_ (.A(_05892_),
    .X(_07526_));
 sky130_fd_sc_hd__a211o_1 _24302_ (.A1(_05527_),
    .A2(_07494_),
    .B1(_07526_),
    .C1(_07503_),
    .X(_07527_));
 sky130_fd_sc_hd__nand2_1 _24303_ (.A(_07498_),
    .B(net1492),
    .Y(_07528_));
 sky130_fd_sc_hd__o21ai_1 _24304_ (.A1(_07521_),
    .A2(_07527_),
    .B1(net1493),
    .Y(_02149_));
 sky130_fd_sc_hd__a211o_1 _24305_ (.A1(_05530_),
    .A2(_07494_),
    .B1(_07526_),
    .C1(_07506_),
    .X(_07529_));
 sky130_fd_sc_hd__nand2_1 _24306_ (.A(_07498_),
    .B(net464),
    .Y(_07530_));
 sky130_fd_sc_hd__o21ai_1 _24307_ (.A1(_07521_),
    .A2(_07529_),
    .B1(net465),
    .Y(_02150_));
 sky130_fd_sc_hd__a211o_1 _24308_ (.A1(_05533_),
    .A2(_07494_),
    .B1(_07526_),
    .C1(_07509_),
    .X(_07531_));
 sky130_fd_sc_hd__nand2_1 _24309_ (.A(_07498_),
    .B(net432),
    .Y(_07532_));
 sky130_fd_sc_hd__o21ai_1 _24310_ (.A1(_07521_),
    .A2(_07531_),
    .B1(net433),
    .Y(_02151_));
 sky130_fd_sc_hd__a211o_1 _24311_ (.A1(_05536_),
    .A2(_07494_),
    .B1(_07526_),
    .C1(_07512_),
    .X(_07533_));
 sky130_fd_sc_hd__nand2_1 _24312_ (.A(_07498_),
    .B(net1144),
    .Y(_07534_));
 sky130_fd_sc_hd__o21ai_1 _24313_ (.A1(_07521_),
    .A2(_07533_),
    .B1(net1145),
    .Y(_02152_));
 sky130_fd_sc_hd__a211o_1 _24314_ (.A1(_05539_),
    .A2(_07494_),
    .B1(_07526_),
    .C1(_07515_),
    .X(_07535_));
 sky130_fd_sc_hd__nand2_1 _24315_ (.A(_07498_),
    .B(net1750),
    .Y(_07536_));
 sky130_fd_sc_hd__o21ai_1 _24316_ (.A1(_07521_),
    .A2(_07535_),
    .B1(net1751),
    .Y(_02153_));
 sky130_fd_sc_hd__a211o_1 _24317_ (.A1(_05542_),
    .A2(_07494_),
    .B1(_07526_),
    .C1(_07518_),
    .X(_07537_));
 sky130_fd_sc_hd__nand2_1 _24318_ (.A(_07498_),
    .B(net1692),
    .Y(_07538_));
 sky130_fd_sc_hd__o21ai_1 _24319_ (.A1(_07521_),
    .A2(_07537_),
    .B1(net1693),
    .Y(_02154_));
 sky130_fd_sc_hd__a211o_1 _24320_ (.A1(_05545_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07496_),
    .X(_07539_));
 sky130_fd_sc_hd__nand2_1 _24321_ (.A(_07493_),
    .B(net1256),
    .Y(_07540_));
 sky130_fd_sc_hd__o21ai_1 _24322_ (.A1(_07521_),
    .A2(_07539_),
    .B1(net1257),
    .Y(_02155_));
 sky130_fd_sc_hd__a211o_1 _24323_ (.A1(_05548_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07500_),
    .X(_07541_));
 sky130_fd_sc_hd__nand2_1 _24324_ (.A(_07493_),
    .B(net1770),
    .Y(_07542_));
 sky130_fd_sc_hd__o21ai_1 _24325_ (.A1(_07521_),
    .A2(_07541_),
    .B1(net1771),
    .Y(_02156_));
 sky130_fd_sc_hd__a211o_1 _24326_ (.A1(_05551_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07503_),
    .X(_07543_));
 sky130_fd_sc_hd__nand2_1 _24327_ (.A(_07493_),
    .B(net1738),
    .Y(_07544_));
 sky130_fd_sc_hd__o21ai_1 _24328_ (.A1(_07521_),
    .A2(_07543_),
    .B1(net1739),
    .Y(_02157_));
 sky130_fd_sc_hd__a211o_1 _24329_ (.A1(_05555_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07506_),
    .X(_07545_));
 sky130_fd_sc_hd__nand2_1 _24330_ (.A(_07493_),
    .B(net1784),
    .Y(_07546_));
 sky130_fd_sc_hd__o21ai_1 _24331_ (.A1(_07521_),
    .A2(_07545_),
    .B1(net1785),
    .Y(_02158_));
 sky130_fd_sc_hd__a211o_1 _24332_ (.A1(_05558_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07509_),
    .X(_07547_));
 sky130_fd_sc_hd__nand2_1 _24333_ (.A(_07493_),
    .B(net1464),
    .Y(_07548_));
 sky130_fd_sc_hd__o21ai_1 _24334_ (.A1(_07521_),
    .A2(_07547_),
    .B1(net1465),
    .Y(_02159_));
 sky130_fd_sc_hd__a211o_1 _24335_ (.A1(_05561_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07512_),
    .X(_07549_));
 sky130_fd_sc_hd__nand2_1 _24336_ (.A(_07493_),
    .B(net1152),
    .Y(_07550_));
 sky130_fd_sc_hd__o21ai_1 _24337_ (.A1(_07521_),
    .A2(_07549_),
    .B1(net1153),
    .Y(_02160_));
 sky130_fd_sc_hd__a211o_1 _24338_ (.A1(_05564_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07515_),
    .X(_07551_));
 sky130_fd_sc_hd__nand2_1 _24339_ (.A(_07493_),
    .B(net1905),
    .Y(_07552_));
 sky130_fd_sc_hd__o21ai_1 _24340_ (.A1(_07521_),
    .A2(_07551_),
    .B1(net1906),
    .Y(_02161_));
 sky130_fd_sc_hd__a211o_1 _24341_ (.A1(_05567_),
    .A2(_07495_),
    .B1(_07526_),
    .C1(_07518_),
    .X(_07553_));
 sky130_fd_sc_hd__nand2_1 _24342_ (.A(_07493_),
    .B(net1989),
    .Y(_07554_));
 sky130_fd_sc_hd__o21ai_1 _24343_ (.A1(_07521_),
    .A2(_07553_),
    .B1(_07554_),
    .Y(_02162_));
 sky130_fd_sc_hd__nand2_1 _24344_ (.A(_04257_),
    .B(_12311_),
    .Y(_07555_));
 sky130_fd_sc_hd__inv_2 _24345_ (.A(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__o21ai_4 _24346_ (.A1(_06755_),
    .A2(_07556_),
    .B1(_06020_),
    .Y(_07557_));
 sky130_fd_sc_hd__mux2_1 _24347_ (.A0(_06530_),
    .A1(net3172),
    .S(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__clkbuf_1 _24348_ (.A(_07558_),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _24349_ (.A0(_06538_),
    .A1(net3356),
    .S(_07557_),
    .X(_07559_));
 sky130_fd_sc_hd__clkbuf_1 _24350_ (.A(_07559_),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _24351_ (.A0(_06540_),
    .A1(net3348),
    .S(_07557_),
    .X(_07560_));
 sky130_fd_sc_hd__clkbuf_1 _24352_ (.A(_07560_),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _24353_ (.A0(_06542_),
    .A1(net3077),
    .S(_07557_),
    .X(_07561_));
 sky130_fd_sc_hd__clkbuf_1 _24354_ (.A(_07561_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _24355_ (.A0(_06544_),
    .A1(net2917),
    .S(_07557_),
    .X(_07562_));
 sky130_fd_sc_hd__clkbuf_1 _24356_ (.A(_07562_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_1 _24357_ (.A0(_06546_),
    .A1(net3397),
    .S(_07557_),
    .X(_07563_));
 sky130_fd_sc_hd__clkbuf_1 _24358_ (.A(_07563_),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _24359_ (.A0(_06548_),
    .A1(net3536),
    .S(_07557_),
    .X(_07564_));
 sky130_fd_sc_hd__clkbuf_1 _24360_ (.A(_07564_),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _24361_ (.A0(_06550_),
    .A1(net2403),
    .S(_07557_),
    .X(_07565_));
 sky130_fd_sc_hd__clkbuf_1 _24362_ (.A(_07565_),
    .X(_02170_));
 sky130_fd_sc_hd__buf_4 _24363_ (.A(_07557_),
    .X(_07566_));
 sky130_fd_sc_hd__buf_4 _24364_ (.A(_07556_),
    .X(_07567_));
 sky130_fd_sc_hd__buf_4 _24365_ (.A(_07556_),
    .X(_07568_));
 sky130_fd_sc_hd__nor2_1 _24366_ (.A(_05583_),
    .B(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__a211o_1 _24367_ (.A1(_05484_),
    .A2(_07567_),
    .B1(_07526_),
    .C1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__buf_4 _24368_ (.A(_07557_),
    .X(_07571_));
 sky130_fd_sc_hd__nand2_1 _24369_ (.A(_07571_),
    .B(net768),
    .Y(_07572_));
 sky130_fd_sc_hd__o21ai_1 _24370_ (.A1(_07566_),
    .A2(_07570_),
    .B1(net769),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _24371_ (.A(_05589_),
    .B(_07568_),
    .Y(_07573_));
 sky130_fd_sc_hd__a211o_1 _24372_ (.A1(_05491_),
    .A2(_07567_),
    .B1(_07526_),
    .C1(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__nand2_1 _24373_ (.A(_07571_),
    .B(net934),
    .Y(_07575_));
 sky130_fd_sc_hd__o21ai_1 _24374_ (.A1(_07566_),
    .A2(_07574_),
    .B1(net935),
    .Y(_02172_));
 sky130_fd_sc_hd__buf_4 _24375_ (.A(_05892_),
    .X(_07576_));
 sky130_fd_sc_hd__nor2_1 _24376_ (.A(_05593_),
    .B(_07568_),
    .Y(_07577_));
 sky130_fd_sc_hd__a211o_1 _24377_ (.A1(_05495_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__nand2_1 _24378_ (.A(_07571_),
    .B(net1836),
    .Y(_07579_));
 sky130_fd_sc_hd__o21ai_1 _24379_ (.A1(_07566_),
    .A2(_07578_),
    .B1(net1837),
    .Y(_02173_));
 sky130_fd_sc_hd__nor2_1 _24380_ (.A(_05597_),
    .B(_07568_),
    .Y(_07580_));
 sky130_fd_sc_hd__a211o_1 _24381_ (.A1(_05500_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07580_),
    .X(_07581_));
 sky130_fd_sc_hd__nand2_1 _24382_ (.A(_07571_),
    .B(net1778),
    .Y(_07582_));
 sky130_fd_sc_hd__o21ai_1 _24383_ (.A1(_07566_),
    .A2(_07581_),
    .B1(net1779),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _24384_ (.A(_05601_),
    .B(_07568_),
    .Y(_07583_));
 sky130_fd_sc_hd__a211o_1 _24385_ (.A1(_05504_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07583_),
    .X(_07584_));
 sky130_fd_sc_hd__nand2_1 _24386_ (.A(_07571_),
    .B(net1732),
    .Y(_07585_));
 sky130_fd_sc_hd__o21ai_1 _24387_ (.A1(_07566_),
    .A2(_07584_),
    .B1(net1733),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _24388_ (.A(_05605_),
    .B(_07568_),
    .Y(_07586_));
 sky130_fd_sc_hd__a211o_1 _24389_ (.A1(_05508_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__nand2_1 _24390_ (.A(_07571_),
    .B(net1640),
    .Y(_07588_));
 sky130_fd_sc_hd__o21ai_1 _24391_ (.A1(_07566_),
    .A2(_07587_),
    .B1(net1641),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _24392_ (.A(_05609_),
    .B(_07568_),
    .Y(_07589_));
 sky130_fd_sc_hd__a211o_1 _24393_ (.A1(_05512_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__nand2_1 _24394_ (.A(_07571_),
    .B(net862),
    .Y(_07591_));
 sky130_fd_sc_hd__o21ai_1 _24395_ (.A1(_07566_),
    .A2(_07590_),
    .B1(net863),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _24396_ (.A(_05613_),
    .B(_07568_),
    .Y(_07592_));
 sky130_fd_sc_hd__a211o_1 _24397_ (.A1(_05516_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__nand2_1 _24398_ (.A(_07571_),
    .B(net1132),
    .Y(_07594_));
 sky130_fd_sc_hd__o21ai_1 _24399_ (.A1(_07566_),
    .A2(_07593_),
    .B1(net1133),
    .Y(_02178_));
 sky130_fd_sc_hd__buf_4 _24400_ (.A(_07557_),
    .X(_07595_));
 sky130_fd_sc_hd__a211o_1 _24401_ (.A1(_05521_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07569_),
    .X(_07596_));
 sky130_fd_sc_hd__nand2_1 _24402_ (.A(_07571_),
    .B(net808),
    .Y(_07597_));
 sky130_fd_sc_hd__o21ai_1 _24403_ (.A1(_07595_),
    .A2(_07596_),
    .B1(net809),
    .Y(_02179_));
 sky130_fd_sc_hd__a211o_1 _24404_ (.A1(_05524_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07573_),
    .X(_07598_));
 sky130_fd_sc_hd__nand2_1 _24405_ (.A(_07571_),
    .B(net742),
    .Y(_07599_));
 sky130_fd_sc_hd__o21ai_1 _24406_ (.A1(_07595_),
    .A2(_07598_),
    .B1(net743),
    .Y(_02180_));
 sky130_fd_sc_hd__a211o_1 _24407_ (.A1(_05527_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07577_),
    .X(_07600_));
 sky130_fd_sc_hd__nand2_1 _24408_ (.A(_07571_),
    .B(net1574),
    .Y(_07601_));
 sky130_fd_sc_hd__o21ai_1 _24409_ (.A1(_07595_),
    .A2(_07600_),
    .B1(net1575),
    .Y(_02181_));
 sky130_fd_sc_hd__a211o_1 _24410_ (.A1(_05530_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07580_),
    .X(_07602_));
 sky130_fd_sc_hd__nand2_1 _24411_ (.A(_07571_),
    .B(net1946),
    .Y(_07603_));
 sky130_fd_sc_hd__o21ai_1 _24412_ (.A1(_07595_),
    .A2(_07602_),
    .B1(net1947),
    .Y(_02182_));
 sky130_fd_sc_hd__a211o_1 _24413_ (.A1(_05533_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07583_),
    .X(_07604_));
 sky130_fd_sc_hd__nand2_1 _24414_ (.A(_07571_),
    .B(net944),
    .Y(_07605_));
 sky130_fd_sc_hd__o21ai_1 _24415_ (.A1(_07595_),
    .A2(_07604_),
    .B1(net945),
    .Y(_02183_));
 sky130_fd_sc_hd__a211o_1 _24416_ (.A1(_05536_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07586_),
    .X(_07606_));
 sky130_fd_sc_hd__nand2_1 _24417_ (.A(_07571_),
    .B(net1258),
    .Y(_07607_));
 sky130_fd_sc_hd__o21ai_1 _24418_ (.A1(_07595_),
    .A2(_07606_),
    .B1(net1259),
    .Y(_02184_));
 sky130_fd_sc_hd__a211o_1 _24419_ (.A1(_05539_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07589_),
    .X(_07608_));
 sky130_fd_sc_hd__nand2_1 _24420_ (.A(_07571_),
    .B(net1476),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_1 _24421_ (.A1(_07595_),
    .A2(_07608_),
    .B1(net1477),
    .Y(_02185_));
 sky130_fd_sc_hd__a211o_1 _24422_ (.A1(_05542_),
    .A2(_07567_),
    .B1(_07576_),
    .C1(_07592_),
    .X(_07610_));
 sky130_fd_sc_hd__nand2_1 _24423_ (.A(_07571_),
    .B(net1706),
    .Y(_07611_));
 sky130_fd_sc_hd__o21ai_1 _24424_ (.A1(_07595_),
    .A2(_07610_),
    .B1(net1707),
    .Y(_02186_));
 sky130_fd_sc_hd__a211o_1 _24425_ (.A1(_05545_),
    .A2(_07568_),
    .B1(_07576_),
    .C1(_07569_),
    .X(_07612_));
 sky130_fd_sc_hd__nand2_1 _24426_ (.A(_07566_),
    .B(net1913),
    .Y(_07613_));
 sky130_fd_sc_hd__o21ai_1 _24427_ (.A1(_07595_),
    .A2(_07612_),
    .B1(net1914),
    .Y(_02187_));
 sky130_fd_sc_hd__a211o_1 _24428_ (.A1(_05548_),
    .A2(_07568_),
    .B1(_07576_),
    .C1(_07573_),
    .X(_07614_));
 sky130_fd_sc_hd__nand2_1 _24429_ (.A(_07566_),
    .B(net1854),
    .Y(_07615_));
 sky130_fd_sc_hd__o21ai_1 _24430_ (.A1(_07595_),
    .A2(_07614_),
    .B1(net1855),
    .Y(_02188_));
 sky130_fd_sc_hd__buf_4 _24431_ (.A(_09057_),
    .X(_07616_));
 sky130_fd_sc_hd__a211o_1 _24432_ (.A1(_05551_),
    .A2(_07568_),
    .B1(_07616_),
    .C1(_07577_),
    .X(_07617_));
 sky130_fd_sc_hd__nand2_1 _24433_ (.A(_07566_),
    .B(net1921),
    .Y(_07618_));
 sky130_fd_sc_hd__o21ai_1 _24434_ (.A1(_07595_),
    .A2(_07617_),
    .B1(net1922),
    .Y(_02189_));
 sky130_fd_sc_hd__a211o_1 _24435_ (.A1(_05555_),
    .A2(_07568_),
    .B1(_07616_),
    .C1(_07580_),
    .X(_07619_));
 sky130_fd_sc_hd__nand2_1 _24436_ (.A(_07566_),
    .B(net1988),
    .Y(_07620_));
 sky130_fd_sc_hd__o21ai_1 _24437_ (.A1(_07595_),
    .A2(_07619_),
    .B1(_07620_),
    .Y(_02190_));
 sky130_fd_sc_hd__a211o_1 _24438_ (.A1(_05558_),
    .A2(_07568_),
    .B1(_07616_),
    .C1(_07583_),
    .X(_07621_));
 sky130_fd_sc_hd__nand2_1 _24439_ (.A(_07566_),
    .B(net1991),
    .Y(_07622_));
 sky130_fd_sc_hd__o21ai_1 _24440_ (.A1(_07595_),
    .A2(_07621_),
    .B1(_07622_),
    .Y(_02191_));
 sky130_fd_sc_hd__a211o_1 _24441_ (.A1(_05561_),
    .A2(_07568_),
    .B1(_07616_),
    .C1(_07586_),
    .X(_07623_));
 sky130_fd_sc_hd__nand2_1 _24442_ (.A(_07566_),
    .B(net1903),
    .Y(_07624_));
 sky130_fd_sc_hd__o21ai_1 _24443_ (.A1(_07595_),
    .A2(_07623_),
    .B1(net1904),
    .Y(_02192_));
 sky130_fd_sc_hd__a211o_1 _24444_ (.A1(_05564_),
    .A2(_07568_),
    .B1(_07616_),
    .C1(_07589_),
    .X(_07625_));
 sky130_fd_sc_hd__nand2_1 _24445_ (.A(_07566_),
    .B(net1867),
    .Y(_07626_));
 sky130_fd_sc_hd__o21ai_1 _24446_ (.A1(_07595_),
    .A2(_07625_),
    .B1(net1868),
    .Y(_02193_));
 sky130_fd_sc_hd__a211o_1 _24447_ (.A1(_05567_),
    .A2(_07568_),
    .B1(_07616_),
    .C1(_07592_),
    .X(_07627_));
 sky130_fd_sc_hd__nand2_1 _24448_ (.A(_07566_),
    .B(net1698),
    .Y(_07628_));
 sky130_fd_sc_hd__o21ai_1 _24449_ (.A1(_07595_),
    .A2(_07627_),
    .B1(net1699),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_4 _24450_ (.A(_12309_),
    .B(_09071_),
    .Y(_07629_));
 sky130_fd_sc_hd__inv_2 _24451_ (.A(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__o21ai_2 _24452_ (.A1(_12289_),
    .A2(_07630_),
    .B1(_12190_),
    .Y(_07631_));
 sky130_fd_sc_hd__clkbuf_8 _24453_ (.A(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__mux2_1 _24454_ (.A0(_06530_),
    .A1(net2504),
    .S(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__clkbuf_1 _24455_ (.A(_07633_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _24456_ (.A0(_06538_),
    .A1(net2363),
    .S(_07632_),
    .X(_07634_));
 sky130_fd_sc_hd__clkbuf_1 _24457_ (.A(_07634_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _24458_ (.A0(_06540_),
    .A1(net2641),
    .S(_07632_),
    .X(_07635_));
 sky130_fd_sc_hd__clkbuf_1 _24459_ (.A(_07635_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _24460_ (.A0(_06542_),
    .A1(net3054),
    .S(_07632_),
    .X(_07636_));
 sky130_fd_sc_hd__clkbuf_1 _24461_ (.A(_07636_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _24462_ (.A0(_06544_),
    .A1(net2251),
    .S(_07632_),
    .X(_07637_));
 sky130_fd_sc_hd__clkbuf_1 _24463_ (.A(_07637_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _24464_ (.A0(_06546_),
    .A1(net3605),
    .S(_07632_),
    .X(_07638_));
 sky130_fd_sc_hd__clkbuf_1 _24465_ (.A(_07638_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _24466_ (.A0(_06548_),
    .A1(net2936),
    .S(_07632_),
    .X(_07639_));
 sky130_fd_sc_hd__clkbuf_1 _24467_ (.A(_07639_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _24468_ (.A0(_06550_),
    .A1(net2949),
    .S(_07632_),
    .X(_07640_));
 sky130_fd_sc_hd__clkbuf_1 _24469_ (.A(_07640_),
    .X(_02202_));
 sky130_fd_sc_hd__buf_4 _24470_ (.A(_07630_),
    .X(_07641_));
 sky130_fd_sc_hd__a21o_1 _24471_ (.A1(_07629_),
    .A2(_12184_),
    .B1(_12851_),
    .X(_07642_));
 sky130_fd_sc_hd__a21oi_1 _24472_ (.A1(_02852_),
    .A2(_07641_),
    .B1(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__mux2_1 _24473_ (.A0(_07643_),
    .A1(net2959),
    .S(_07632_),
    .X(_07644_));
 sky130_fd_sc_hd__clkbuf_1 _24474_ (.A(_07644_),
    .X(_02203_));
 sky130_fd_sc_hd__a21o_1 _24475_ (.A1(_07629_),
    .A2(_12197_),
    .B1(_12851_),
    .X(_07645_));
 sky130_fd_sc_hd__a21oi_1 _24476_ (.A1(_02862_),
    .A2(_07641_),
    .B1(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__mux2_1 _24477_ (.A0(_07646_),
    .A1(net3507),
    .S(_07632_),
    .X(_07647_));
 sky130_fd_sc_hd__clkbuf_1 _24478_ (.A(_07647_),
    .X(_02204_));
 sky130_fd_sc_hd__a21o_1 _24479_ (.A1(_07629_),
    .A2(_12205_),
    .B1(_12851_),
    .X(_07648_));
 sky130_fd_sc_hd__a21oi_1 _24480_ (.A1(_02869_),
    .A2(_07641_),
    .B1(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__mux2_1 _24481_ (.A0(_07649_),
    .A1(net3699),
    .S(_07632_),
    .X(_07650_));
 sky130_fd_sc_hd__clkbuf_1 _24482_ (.A(_07650_),
    .X(_02205_));
 sky130_fd_sc_hd__a21o_1 _24483_ (.A1(_07629_),
    .A2(_12213_),
    .B1(_12851_),
    .X(_07651_));
 sky130_fd_sc_hd__a21oi_1 _24484_ (.A1(_02876_),
    .A2(_07641_),
    .B1(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__mux2_1 _24485_ (.A0(_07652_),
    .A1(net3659),
    .S(_07632_),
    .X(_07653_));
 sky130_fd_sc_hd__clkbuf_1 _24486_ (.A(_07653_),
    .X(_02206_));
 sky130_fd_sc_hd__a21o_1 _24487_ (.A1(_07629_),
    .A2(_12221_),
    .B1(_12851_),
    .X(_07654_));
 sky130_fd_sc_hd__a21oi_1 _24488_ (.A1(_02883_),
    .A2(_07641_),
    .B1(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__mux2_1 _24489_ (.A0(_07655_),
    .A1(net3647),
    .S(_07632_),
    .X(_07656_));
 sky130_fd_sc_hd__clkbuf_1 _24490_ (.A(_07656_),
    .X(_02207_));
 sky130_fd_sc_hd__a21o_1 _24491_ (.A1(_07629_),
    .A2(_12229_),
    .B1(_09129_),
    .X(_07657_));
 sky130_fd_sc_hd__a21oi_1 _24492_ (.A1(_02890_),
    .A2(_07641_),
    .B1(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__mux2_1 _24493_ (.A0(_07658_),
    .A1(net3766),
    .S(_07632_),
    .X(_07659_));
 sky130_fd_sc_hd__clkbuf_1 _24494_ (.A(_07659_),
    .X(_02208_));
 sky130_fd_sc_hd__a21o_1 _24495_ (.A1(_07629_),
    .A2(_12237_),
    .B1(_09129_),
    .X(_07660_));
 sky130_fd_sc_hd__a21oi_1 _24496_ (.A1(_02897_),
    .A2(_07641_),
    .B1(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__mux2_1 _24497_ (.A0(_07661_),
    .A1(net3586),
    .S(_07632_),
    .X(_07662_));
 sky130_fd_sc_hd__clkbuf_1 _24498_ (.A(_07662_),
    .X(_02209_));
 sky130_fd_sc_hd__a21o_1 _24499_ (.A1(_07629_),
    .A2(_12245_),
    .B1(_09129_),
    .X(_07663_));
 sky130_fd_sc_hd__a21oi_1 _24500_ (.A1(_02904_),
    .A2(_07641_),
    .B1(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__mux2_1 _24501_ (.A0(_07664_),
    .A1(net3312),
    .S(_07632_),
    .X(_07665_));
 sky130_fd_sc_hd__clkbuf_1 _24502_ (.A(_07665_),
    .X(_02210_));
 sky130_fd_sc_hd__a21oi_1 _24503_ (.A1(_02912_),
    .A2(_07641_),
    .B1(_07642_),
    .Y(_07666_));
 sky130_fd_sc_hd__buf_6 _24504_ (.A(_07631_),
    .X(_07667_));
 sky130_fd_sc_hd__mux2_1 _24505_ (.A0(_07666_),
    .A1(net3159),
    .S(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__clkbuf_1 _24506_ (.A(_07668_),
    .X(_02211_));
 sky130_fd_sc_hd__a21oi_1 _24507_ (.A1(_02917_),
    .A2(_07641_),
    .B1(_07645_),
    .Y(_07669_));
 sky130_fd_sc_hd__mux2_1 _24508_ (.A0(_07669_),
    .A1(net3380),
    .S(_07667_),
    .X(_07670_));
 sky130_fd_sc_hd__clkbuf_1 _24509_ (.A(_07670_),
    .X(_02212_));
 sky130_fd_sc_hd__a21oi_1 _24510_ (.A1(_02922_),
    .A2(_07641_),
    .B1(_07648_),
    .Y(_07671_));
 sky130_fd_sc_hd__mux2_1 _24511_ (.A0(_07671_),
    .A1(net3250),
    .S(_07667_),
    .X(_07672_));
 sky130_fd_sc_hd__clkbuf_1 _24512_ (.A(_07672_),
    .X(_02213_));
 sky130_fd_sc_hd__a21oi_1 _24513_ (.A1(_02928_),
    .A2(_07641_),
    .B1(_07651_),
    .Y(_07673_));
 sky130_fd_sc_hd__mux2_1 _24514_ (.A0(_07673_),
    .A1(net3794),
    .S(_07667_),
    .X(_07674_));
 sky130_fd_sc_hd__clkbuf_1 _24515_ (.A(_07674_),
    .X(_02214_));
 sky130_fd_sc_hd__a21oi_1 _24516_ (.A1(_02933_),
    .A2(_07641_),
    .B1(_07654_),
    .Y(_07675_));
 sky130_fd_sc_hd__mux2_1 _24517_ (.A0(_07675_),
    .A1(net3535),
    .S(_07667_),
    .X(_07676_));
 sky130_fd_sc_hd__clkbuf_1 _24518_ (.A(_07676_),
    .X(_02215_));
 sky130_fd_sc_hd__a21oi_1 _24519_ (.A1(_02938_),
    .A2(_07641_),
    .B1(_07657_),
    .Y(_07677_));
 sky130_fd_sc_hd__mux2_1 _24520_ (.A0(_07677_),
    .A1(net3748),
    .S(_07667_),
    .X(_07678_));
 sky130_fd_sc_hd__clkbuf_1 _24521_ (.A(_07678_),
    .X(_02216_));
 sky130_fd_sc_hd__a21oi_1 _24522_ (.A1(_02943_),
    .A2(_07641_),
    .B1(_07660_),
    .Y(_07679_));
 sky130_fd_sc_hd__mux2_1 _24523_ (.A0(_07679_),
    .A1(net3693),
    .S(_07667_),
    .X(_07680_));
 sky130_fd_sc_hd__clkbuf_1 _24524_ (.A(_07680_),
    .X(_02217_));
 sky130_fd_sc_hd__a21oi_1 _24525_ (.A1(_02948_),
    .A2(_07641_),
    .B1(_07663_),
    .Y(_07681_));
 sky130_fd_sc_hd__mux2_1 _24526_ (.A0(_07681_),
    .A1(net3262),
    .S(_07667_),
    .X(_07682_));
 sky130_fd_sc_hd__clkbuf_1 _24527_ (.A(_07682_),
    .X(_02218_));
 sky130_fd_sc_hd__a21oi_1 _24528_ (.A1(_02952_),
    .A2(_07630_),
    .B1(_07642_),
    .Y(_07683_));
 sky130_fd_sc_hd__mux2_1 _24529_ (.A0(_07683_),
    .A1(net3933),
    .S(_07667_),
    .X(_07684_));
 sky130_fd_sc_hd__clkbuf_1 _24530_ (.A(_07684_),
    .X(_02219_));
 sky130_fd_sc_hd__a21oi_1 _24531_ (.A1(_02956_),
    .A2(_07630_),
    .B1(_07645_),
    .Y(_07685_));
 sky130_fd_sc_hd__mux2_1 _24532_ (.A0(_07685_),
    .A1(net3673),
    .S(_07667_),
    .X(_07686_));
 sky130_fd_sc_hd__clkbuf_1 _24533_ (.A(_07686_),
    .X(_02220_));
 sky130_fd_sc_hd__a21oi_1 _24534_ (.A1(_02960_),
    .A2(_07630_),
    .B1(_07648_),
    .Y(_07687_));
 sky130_fd_sc_hd__mux2_1 _24535_ (.A0(_07687_),
    .A1(net3807),
    .S(_07667_),
    .X(_07688_));
 sky130_fd_sc_hd__clkbuf_1 _24536_ (.A(_07688_),
    .X(_02221_));
 sky130_fd_sc_hd__a21oi_1 _24537_ (.A1(_02964_),
    .A2(_07630_),
    .B1(_07651_),
    .Y(_07689_));
 sky130_fd_sc_hd__mux2_1 _24538_ (.A0(_07689_),
    .A1(net3671),
    .S(_07667_),
    .X(_07690_));
 sky130_fd_sc_hd__clkbuf_1 _24539_ (.A(_07690_),
    .X(_02222_));
 sky130_fd_sc_hd__a21oi_1 _24540_ (.A1(_02968_),
    .A2(_07630_),
    .B1(_07654_),
    .Y(_07691_));
 sky130_fd_sc_hd__mux2_1 _24541_ (.A0(_07691_),
    .A1(net3779),
    .S(_07667_),
    .X(_07692_));
 sky130_fd_sc_hd__clkbuf_1 _24542_ (.A(_07692_),
    .X(_02223_));
 sky130_fd_sc_hd__a21oi_1 _24543_ (.A1(_02972_),
    .A2(_07630_),
    .B1(_07657_),
    .Y(_07693_));
 sky130_fd_sc_hd__mux2_1 _24544_ (.A0(_07693_),
    .A1(net3946),
    .S(_07667_),
    .X(_07694_));
 sky130_fd_sc_hd__clkbuf_1 _24545_ (.A(_07694_),
    .X(_02224_));
 sky130_fd_sc_hd__a21oi_1 _24546_ (.A1(_02976_),
    .A2(_07630_),
    .B1(_07660_),
    .Y(_07695_));
 sky130_fd_sc_hd__mux2_1 _24547_ (.A0(_07695_),
    .A1(net3955),
    .S(_07667_),
    .X(_07696_));
 sky130_fd_sc_hd__clkbuf_1 _24548_ (.A(_07696_),
    .X(_02225_));
 sky130_fd_sc_hd__a21oi_1 _24549_ (.A1(_02980_),
    .A2(_07630_),
    .B1(_07663_),
    .Y(_07697_));
 sky130_fd_sc_hd__mux2_1 _24550_ (.A0(_07697_),
    .A1(net3941),
    .S(_07667_),
    .X(_07698_));
 sky130_fd_sc_hd__clkbuf_1 _24551_ (.A(_07698_),
    .X(_02226_));
 sky130_fd_sc_hd__buf_6 _24552_ (.A(_02809_),
    .X(_07699_));
 sky130_fd_sc_hd__nor2_2 _24553_ (.A(_12313_),
    .B(_02816_),
    .Y(_07700_));
 sky130_fd_sc_hd__o21ai_4 _24554_ (.A1(_06755_),
    .A2(_07700_),
    .B1(_12190_),
    .Y(_07701_));
 sky130_fd_sc_hd__mux2_1 _24555_ (.A0(_07699_),
    .A1(net2284),
    .S(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__clkbuf_1 _24556_ (.A(_07702_),
    .X(_02227_));
 sky130_fd_sc_hd__buf_8 _24557_ (.A(_02822_),
    .X(_07703_));
 sky130_fd_sc_hd__mux2_1 _24558_ (.A0(_07703_),
    .A1(net2344),
    .S(_07701_),
    .X(_07704_));
 sky130_fd_sc_hd__clkbuf_1 _24559_ (.A(_07704_),
    .X(_02228_));
 sky130_fd_sc_hd__buf_8 _24560_ (.A(_02826_),
    .X(_07705_));
 sky130_fd_sc_hd__mux2_1 _24561_ (.A0(_07705_),
    .A1(net2040),
    .S(_07701_),
    .X(_07706_));
 sky130_fd_sc_hd__clkbuf_1 _24562_ (.A(_07706_),
    .X(_02229_));
 sky130_fd_sc_hd__buf_8 _24563_ (.A(_02830_),
    .X(_07707_));
 sky130_fd_sc_hd__mux2_1 _24564_ (.A0(_07707_),
    .A1(net2210),
    .S(_07701_),
    .X(_07708_));
 sky130_fd_sc_hd__clkbuf_1 _24565_ (.A(_07708_),
    .X(_02230_));
 sky130_fd_sc_hd__buf_8 _24566_ (.A(_02834_),
    .X(_07709_));
 sky130_fd_sc_hd__mux2_1 _24567_ (.A0(_07709_),
    .A1(net3152),
    .S(_07701_),
    .X(_07710_));
 sky130_fd_sc_hd__clkbuf_1 _24568_ (.A(_07710_),
    .X(_02231_));
 sky130_fd_sc_hd__buf_8 _24569_ (.A(_02838_),
    .X(_07711_));
 sky130_fd_sc_hd__mux2_1 _24570_ (.A0(_07711_),
    .A1(net2211),
    .S(_07701_),
    .X(_07712_));
 sky130_fd_sc_hd__clkbuf_1 _24571_ (.A(_07712_),
    .X(_02232_));
 sky130_fd_sc_hd__buf_8 _24572_ (.A(_02842_),
    .X(_07713_));
 sky130_fd_sc_hd__mux2_1 _24573_ (.A0(_07713_),
    .A1(net2144),
    .S(_07701_),
    .X(_07714_));
 sky130_fd_sc_hd__clkbuf_1 _24574_ (.A(_07714_),
    .X(_02233_));
 sky130_fd_sc_hd__buf_6 _24575_ (.A(_02846_),
    .X(_07715_));
 sky130_fd_sc_hd__mux2_1 _24576_ (.A0(_07715_),
    .A1(net2103),
    .S(_07701_),
    .X(_07716_));
 sky130_fd_sc_hd__clkbuf_1 _24577_ (.A(_07716_),
    .X(_02234_));
 sky130_fd_sc_hd__buf_4 _24578_ (.A(_07701_),
    .X(_07717_));
 sky130_fd_sc_hd__buf_4 _24579_ (.A(_07700_),
    .X(_07718_));
 sky130_fd_sc_hd__buf_4 _24580_ (.A(_07700_),
    .X(_07719_));
 sky130_fd_sc_hd__nor2_1 _24581_ (.A(_05583_),
    .B(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__a211o_1 _24582_ (.A1(_05484_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__buf_4 _24583_ (.A(_07701_),
    .X(_07722_));
 sky130_fd_sc_hd__nand2_1 _24584_ (.A(_07722_),
    .B(net996),
    .Y(_07723_));
 sky130_fd_sc_hd__o21ai_1 _24585_ (.A1(_07717_),
    .A2(_07721_),
    .B1(net997),
    .Y(_02235_));
 sky130_fd_sc_hd__nor2_1 _24586_ (.A(_05589_),
    .B(_07719_),
    .Y(_07724_));
 sky130_fd_sc_hd__a211o_1 _24587_ (.A1(_05491_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__nand2_1 _24588_ (.A(_07722_),
    .B(net1314),
    .Y(_07726_));
 sky130_fd_sc_hd__o21ai_1 _24589_ (.A1(_07717_),
    .A2(_07725_),
    .B1(net1315),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _24590_ (.A(_05593_),
    .B(_07719_),
    .Y(_07727_));
 sky130_fd_sc_hd__a211o_1 _24591_ (.A1(_05495_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07727_),
    .X(_07728_));
 sky130_fd_sc_hd__nand2_1 _24592_ (.A(_07722_),
    .B(net1644),
    .Y(_07729_));
 sky130_fd_sc_hd__o21ai_1 _24593_ (.A1(_07717_),
    .A2(_07728_),
    .B1(net1645),
    .Y(_02237_));
 sky130_fd_sc_hd__nor2_1 _24594_ (.A(_05597_),
    .B(_07719_),
    .Y(_07730_));
 sky130_fd_sc_hd__a211o_1 _24595_ (.A1(_05500_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__nand2_1 _24596_ (.A(_07722_),
    .B(net394),
    .Y(_07732_));
 sky130_fd_sc_hd__o21ai_1 _24597_ (.A1(_07717_),
    .A2(_07731_),
    .B1(net395),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _24598_ (.A(_05601_),
    .B(_07719_),
    .Y(_07733_));
 sky130_fd_sc_hd__a211o_1 _24599_ (.A1(_05504_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__nand2_1 _24600_ (.A(_07722_),
    .B(net416),
    .Y(_07735_));
 sky130_fd_sc_hd__o21ai_1 _24601_ (.A1(_07717_),
    .A2(_07734_),
    .B1(net417),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _24602_ (.A(_05605_),
    .B(_07719_),
    .Y(_07736_));
 sky130_fd_sc_hd__a211o_1 _24603_ (.A1(_05508_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__nand2_1 _24604_ (.A(_07722_),
    .B(net490),
    .Y(_07738_));
 sky130_fd_sc_hd__o21ai_1 _24605_ (.A1(_07717_),
    .A2(_07737_),
    .B1(net491),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_1 _24606_ (.A(_05609_),
    .B(_07719_),
    .Y(_07739_));
 sky130_fd_sc_hd__a211o_1 _24607_ (.A1(_05512_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__nand2_1 _24608_ (.A(_07722_),
    .B(net1002),
    .Y(_07741_));
 sky130_fd_sc_hd__o21ai_1 _24609_ (.A1(_07717_),
    .A2(_07740_),
    .B1(net1003),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_1 _24610_ (.A(_05613_),
    .B(_07719_),
    .Y(_07742_));
 sky130_fd_sc_hd__a211o_1 _24611_ (.A1(_05516_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__nand2_1 _24612_ (.A(_07722_),
    .B(net558),
    .Y(_07744_));
 sky130_fd_sc_hd__o21ai_1 _24613_ (.A1(_07717_),
    .A2(_07743_),
    .B1(net559),
    .Y(_02242_));
 sky130_fd_sc_hd__buf_4 _24614_ (.A(_07701_),
    .X(_07745_));
 sky130_fd_sc_hd__a211o_1 _24615_ (.A1(_05521_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07720_),
    .X(_07746_));
 sky130_fd_sc_hd__nand2_1 _24616_ (.A(_07722_),
    .B(net1320),
    .Y(_07747_));
 sky130_fd_sc_hd__o21ai_1 _24617_ (.A1(_07745_),
    .A2(_07746_),
    .B1(net1321),
    .Y(_02243_));
 sky130_fd_sc_hd__a211o_1 _24618_ (.A1(_05524_),
    .A2(_07718_),
    .B1(_07616_),
    .C1(_07724_),
    .X(_07748_));
 sky130_fd_sc_hd__nand2_1 _24619_ (.A(_07722_),
    .B(net484),
    .Y(_07749_));
 sky130_fd_sc_hd__o21ai_1 _24620_ (.A1(_07745_),
    .A2(_07748_),
    .B1(net485),
    .Y(_02244_));
 sky130_fd_sc_hd__buf_4 _24621_ (.A(_09057_),
    .X(_07750_));
 sky130_fd_sc_hd__a211o_1 _24622_ (.A1(_05527_),
    .A2(_07718_),
    .B1(_07750_),
    .C1(_07727_),
    .X(_07751_));
 sky130_fd_sc_hd__nand2_1 _24623_ (.A(_07722_),
    .B(net1308),
    .Y(_07752_));
 sky130_fd_sc_hd__o21ai_1 _24624_ (.A1(_07745_),
    .A2(_07751_),
    .B1(net1309),
    .Y(_02245_));
 sky130_fd_sc_hd__a211o_1 _24625_ (.A1(_05530_),
    .A2(_07718_),
    .B1(_07750_),
    .C1(_07730_),
    .X(_07753_));
 sky130_fd_sc_hd__nand2_1 _24626_ (.A(_07722_),
    .B(net448),
    .Y(_07754_));
 sky130_fd_sc_hd__o21ai_1 _24627_ (.A1(_07745_),
    .A2(_07753_),
    .B1(net449),
    .Y(_02246_));
 sky130_fd_sc_hd__a211o_1 _24628_ (.A1(_05533_),
    .A2(_07718_),
    .B1(_07750_),
    .C1(_07733_),
    .X(_07755_));
 sky130_fd_sc_hd__nand2_1 _24629_ (.A(_07722_),
    .B(net1118),
    .Y(_07756_));
 sky130_fd_sc_hd__o21ai_1 _24630_ (.A1(_07745_),
    .A2(_07755_),
    .B1(net1119),
    .Y(_02247_));
 sky130_fd_sc_hd__a211o_1 _24631_ (.A1(_05536_),
    .A2(_07718_),
    .B1(_07750_),
    .C1(_07736_),
    .X(_07757_));
 sky130_fd_sc_hd__nand2_1 _24632_ (.A(_07722_),
    .B(net566),
    .Y(_07758_));
 sky130_fd_sc_hd__o21ai_1 _24633_ (.A1(_07745_),
    .A2(_07757_),
    .B1(net567),
    .Y(_02248_));
 sky130_fd_sc_hd__a211o_1 _24634_ (.A1(_05539_),
    .A2(_07718_),
    .B1(_07750_),
    .C1(_07739_),
    .X(_07759_));
 sky130_fd_sc_hd__nand2_1 _24635_ (.A(_07722_),
    .B(net446),
    .Y(_07760_));
 sky130_fd_sc_hd__o21ai_1 _24636_ (.A1(_07745_),
    .A2(_07759_),
    .B1(net447),
    .Y(_02249_));
 sky130_fd_sc_hd__a211o_1 _24637_ (.A1(_05542_),
    .A2(_07718_),
    .B1(_07750_),
    .C1(_07742_),
    .X(_07761_));
 sky130_fd_sc_hd__nand2_1 _24638_ (.A(_07722_),
    .B(net1790),
    .Y(_07762_));
 sky130_fd_sc_hd__o21ai_1 _24639_ (.A1(_07745_),
    .A2(_07761_),
    .B1(net1791),
    .Y(_02250_));
 sky130_fd_sc_hd__a211o_1 _24640_ (.A1(_05545_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07720_),
    .X(_07763_));
 sky130_fd_sc_hd__nand2_1 _24641_ (.A(_07717_),
    .B(net610),
    .Y(_07764_));
 sky130_fd_sc_hd__o21ai_1 _24642_ (.A1(_07745_),
    .A2(_07763_),
    .B1(net611),
    .Y(_02251_));
 sky130_fd_sc_hd__a211o_1 _24643_ (.A1(_05548_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07724_),
    .X(_07765_));
 sky130_fd_sc_hd__nand2_1 _24644_ (.A(_07717_),
    .B(net454),
    .Y(_07766_));
 sky130_fd_sc_hd__o21ai_1 _24645_ (.A1(_07745_),
    .A2(_07765_),
    .B1(net455),
    .Y(_02252_));
 sky130_fd_sc_hd__a211o_1 _24646_ (.A1(_05551_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07727_),
    .X(_07767_));
 sky130_fd_sc_hd__nand2_1 _24647_ (.A(_07717_),
    .B(net1596),
    .Y(_07768_));
 sky130_fd_sc_hd__o21ai_1 _24648_ (.A1(_07745_),
    .A2(_07767_),
    .B1(net1597),
    .Y(_02253_));
 sky130_fd_sc_hd__a211o_1 _24649_ (.A1(_05555_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07730_),
    .X(_07769_));
 sky130_fd_sc_hd__nand2_1 _24650_ (.A(_07717_),
    .B(net1726),
    .Y(_07770_));
 sky130_fd_sc_hd__o21ai_1 _24651_ (.A1(_07745_),
    .A2(_07769_),
    .B1(net1727),
    .Y(_02254_));
 sky130_fd_sc_hd__a211o_1 _24652_ (.A1(_05558_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07733_),
    .X(_07771_));
 sky130_fd_sc_hd__nand2_1 _24653_ (.A(_07717_),
    .B(net1482),
    .Y(_07772_));
 sky130_fd_sc_hd__o21ai_1 _24654_ (.A1(_07745_),
    .A2(_07771_),
    .B1(net1483),
    .Y(_02255_));
 sky130_fd_sc_hd__a211o_1 _24655_ (.A1(_05561_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07736_),
    .X(_07773_));
 sky130_fd_sc_hd__nand2_1 _24656_ (.A(_07717_),
    .B(net502),
    .Y(_07774_));
 sky130_fd_sc_hd__o21ai_1 _24657_ (.A1(_07745_),
    .A2(_07773_),
    .B1(net503),
    .Y(_02256_));
 sky130_fd_sc_hd__a211o_1 _24658_ (.A1(_05564_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07739_),
    .X(_07775_));
 sky130_fd_sc_hd__nand2_1 _24659_ (.A(_07717_),
    .B(net1332),
    .Y(_07776_));
 sky130_fd_sc_hd__o21ai_1 _24660_ (.A1(_07745_),
    .A2(_07775_),
    .B1(net1333),
    .Y(_02257_));
 sky130_fd_sc_hd__a211o_1 _24661_ (.A1(_05567_),
    .A2(_07719_),
    .B1(_07750_),
    .C1(_07742_),
    .X(_07777_));
 sky130_fd_sc_hd__nand2_1 _24662_ (.A(_07717_),
    .B(net456),
    .Y(_07778_));
 sky130_fd_sc_hd__o21ai_1 _24663_ (.A1(_07745_),
    .A2(_07777_),
    .B1(net457),
    .Y(_02258_));
 sky130_fd_sc_hd__nand2_1 _24664_ (.A(_02983_),
    .B(_12177_),
    .Y(_07779_));
 sky130_fd_sc_hd__inv_2 _24665_ (.A(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__o21ai_4 _24666_ (.A1(_06755_),
    .A2(_07780_),
    .B1(_12190_),
    .Y(_07781_));
 sky130_fd_sc_hd__mux2_1 _24667_ (.A0(_07699_),
    .A1(net2151),
    .S(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__clkbuf_1 _24668_ (.A(_07782_),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _24669_ (.A0(_07703_),
    .A1(net2033),
    .S(_07781_),
    .X(_07783_));
 sky130_fd_sc_hd__clkbuf_1 _24670_ (.A(_07783_),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _24671_ (.A0(_07705_),
    .A1(net2332),
    .S(_07781_),
    .X(_07784_));
 sky130_fd_sc_hd__clkbuf_1 _24672_ (.A(_07784_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _24673_ (.A0(_07707_),
    .A1(net2052),
    .S(_07781_),
    .X(_07785_));
 sky130_fd_sc_hd__clkbuf_1 _24674_ (.A(_07785_),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _24675_ (.A0(_07709_),
    .A1(net2200),
    .S(_07781_),
    .X(_07786_));
 sky130_fd_sc_hd__clkbuf_1 _24676_ (.A(_07786_),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _24677_ (.A0(_07711_),
    .A1(net2916),
    .S(_07781_),
    .X(_07787_));
 sky130_fd_sc_hd__clkbuf_1 _24678_ (.A(_07787_),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _24679_ (.A0(_07713_),
    .A1(net3146),
    .S(_07781_),
    .X(_07788_));
 sky130_fd_sc_hd__clkbuf_1 _24680_ (.A(_07788_),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _24681_ (.A0(_07715_),
    .A1(net3460),
    .S(_07781_),
    .X(_07789_));
 sky130_fd_sc_hd__clkbuf_1 _24682_ (.A(_07789_),
    .X(_02266_));
 sky130_fd_sc_hd__buf_4 _24683_ (.A(_07781_),
    .X(_07790_));
 sky130_fd_sc_hd__buf_4 _24684_ (.A(_07780_),
    .X(_07791_));
 sky130_fd_sc_hd__buf_4 _24685_ (.A(_07780_),
    .X(_07792_));
 sky130_fd_sc_hd__nor2_1 _24686_ (.A(_05583_),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__a211o_1 _24687_ (.A1(_02851_),
    .A2(_07791_),
    .B1(_07750_),
    .C1(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__buf_4 _24688_ (.A(_07781_),
    .X(_07795_));
 sky130_fd_sc_hd__nand2_1 _24689_ (.A(_07795_),
    .B(net562),
    .Y(_07796_));
 sky130_fd_sc_hd__o21ai_1 _24690_ (.A1(_07790_),
    .A2(_07794_),
    .B1(net563),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _24691_ (.A(_05589_),
    .B(_07792_),
    .Y(_07797_));
 sky130_fd_sc_hd__a211o_1 _24692_ (.A1(_02861_),
    .A2(_07791_),
    .B1(_07750_),
    .C1(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__nand2_1 _24693_ (.A(_07795_),
    .B(net1470),
    .Y(_07799_));
 sky130_fd_sc_hd__o21ai_1 _24694_ (.A1(_07790_),
    .A2(_07798_),
    .B1(net1471),
    .Y(_02268_));
 sky130_fd_sc_hd__buf_4 _24695_ (.A(_09057_),
    .X(_07800_));
 sky130_fd_sc_hd__nor2_1 _24696_ (.A(_05593_),
    .B(_07792_),
    .Y(_07801_));
 sky130_fd_sc_hd__a211o_1 _24697_ (.A1(_02868_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__nand2_1 _24698_ (.A(_07795_),
    .B(net1580),
    .Y(_07803_));
 sky130_fd_sc_hd__o21ai_1 _24699_ (.A1(_07790_),
    .A2(_07802_),
    .B1(net1581),
    .Y(_02269_));
 sky130_fd_sc_hd__nor2_1 _24700_ (.A(_05597_),
    .B(_07792_),
    .Y(_07804_));
 sky130_fd_sc_hd__a211o_1 _24701_ (.A1(_02875_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__nand2_1 _24702_ (.A(_07795_),
    .B(net1468),
    .Y(_07806_));
 sky130_fd_sc_hd__o21ai_1 _24703_ (.A1(_07790_),
    .A2(_07805_),
    .B1(net1469),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _24704_ (.A(_05601_),
    .B(_07792_),
    .Y(_07807_));
 sky130_fd_sc_hd__a211o_1 _24705_ (.A1(_02882_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__nand2_1 _24706_ (.A(_07795_),
    .B(net664),
    .Y(_07809_));
 sky130_fd_sc_hd__o21ai_1 _24707_ (.A1(_07790_),
    .A2(_07808_),
    .B1(net665),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _24708_ (.A(_05605_),
    .B(_07792_),
    .Y(_07810_));
 sky130_fd_sc_hd__a211o_1 _24709_ (.A1(_02889_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__nand2_1 _24710_ (.A(_07795_),
    .B(net548),
    .Y(_07812_));
 sky130_fd_sc_hd__o21ai_1 _24711_ (.A1(_07790_),
    .A2(_07811_),
    .B1(net549),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _24712_ (.A(_05609_),
    .B(_07792_),
    .Y(_07813_));
 sky130_fd_sc_hd__a211o_1 _24713_ (.A1(_02896_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__nand2_1 _24714_ (.A(_07795_),
    .B(net1266),
    .Y(_07815_));
 sky130_fd_sc_hd__o21ai_1 _24715_ (.A1(_07790_),
    .A2(_07814_),
    .B1(net1267),
    .Y(_02273_));
 sky130_fd_sc_hd__nor2_1 _24716_ (.A(_05613_),
    .B(_07792_),
    .Y(_07816_));
 sky130_fd_sc_hd__a211o_1 _24717_ (.A1(_02903_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__nand2_1 _24718_ (.A(_07795_),
    .B(net756),
    .Y(_07818_));
 sky130_fd_sc_hd__o21ai_1 _24719_ (.A1(_07790_),
    .A2(_07817_),
    .B1(net757),
    .Y(_02274_));
 sky130_fd_sc_hd__buf_4 _24720_ (.A(_07781_),
    .X(_07819_));
 sky130_fd_sc_hd__a211o_1 _24721_ (.A1(_02911_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07793_),
    .X(_07820_));
 sky130_fd_sc_hd__nand2_1 _24722_ (.A(_07795_),
    .B(net590),
    .Y(_07821_));
 sky130_fd_sc_hd__o21ai_1 _24723_ (.A1(_07819_),
    .A2(_07820_),
    .B1(net591),
    .Y(_02275_));
 sky130_fd_sc_hd__a211o_1 _24724_ (.A1(_02916_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07797_),
    .X(_07822_));
 sky130_fd_sc_hd__nand2_1 _24725_ (.A(_07795_),
    .B(net704),
    .Y(_07823_));
 sky130_fd_sc_hd__o21ai_1 _24726_ (.A1(_07819_),
    .A2(_07822_),
    .B1(net705),
    .Y(_02276_));
 sky130_fd_sc_hd__a211o_1 _24727_ (.A1(_02921_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07801_),
    .X(_07824_));
 sky130_fd_sc_hd__nand2_1 _24728_ (.A(_07795_),
    .B(net1548),
    .Y(_07825_));
 sky130_fd_sc_hd__o21ai_1 _24729_ (.A1(_07819_),
    .A2(_07824_),
    .B1(net1549),
    .Y(_02277_));
 sky130_fd_sc_hd__a211o_1 _24730_ (.A1(_02927_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07804_),
    .X(_07826_));
 sky130_fd_sc_hd__nand2_1 _24731_ (.A(_07795_),
    .B(net696),
    .Y(_07827_));
 sky130_fd_sc_hd__o21ai_1 _24732_ (.A1(_07819_),
    .A2(_07826_),
    .B1(net697),
    .Y(_02278_));
 sky130_fd_sc_hd__a211o_1 _24733_ (.A1(_02932_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07807_),
    .X(_07828_));
 sky130_fd_sc_hd__nand2_1 _24734_ (.A(_07795_),
    .B(net690),
    .Y(_07829_));
 sky130_fd_sc_hd__o21ai_1 _24735_ (.A1(_07819_),
    .A2(_07828_),
    .B1(net691),
    .Y(_02279_));
 sky130_fd_sc_hd__a211o_1 _24736_ (.A1(_02937_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07810_),
    .X(_07830_));
 sky130_fd_sc_hd__nand2_1 _24737_ (.A(_07795_),
    .B(net1016),
    .Y(_07831_));
 sky130_fd_sc_hd__o21ai_1 _24738_ (.A1(_07819_),
    .A2(_07830_),
    .B1(net1017),
    .Y(_02280_));
 sky130_fd_sc_hd__a211o_1 _24739_ (.A1(_02942_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07813_),
    .X(_07832_));
 sky130_fd_sc_hd__nand2_1 _24740_ (.A(_07795_),
    .B(net1356),
    .Y(_07833_));
 sky130_fd_sc_hd__o21ai_1 _24741_ (.A1(_07819_),
    .A2(_07832_),
    .B1(net1357),
    .Y(_02281_));
 sky130_fd_sc_hd__a211o_1 _24742_ (.A1(_02947_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07816_),
    .X(_07834_));
 sky130_fd_sc_hd__nand2_1 _24743_ (.A(_07795_),
    .B(net910),
    .Y(_07835_));
 sky130_fd_sc_hd__o21ai_1 _24744_ (.A1(_07819_),
    .A2(_07834_),
    .B1(net911),
    .Y(_02282_));
 sky130_fd_sc_hd__a211o_1 _24745_ (.A1(_02951_),
    .A2(_07792_),
    .B1(_07800_),
    .C1(_07793_),
    .X(_07836_));
 sky130_fd_sc_hd__nand2_1 _24746_ (.A(_07790_),
    .B(net1388),
    .Y(_07837_));
 sky130_fd_sc_hd__o21ai_1 _24747_ (.A1(_07819_),
    .A2(_07836_),
    .B1(net1389),
    .Y(_02283_));
 sky130_fd_sc_hd__a211o_1 _24748_ (.A1(_02955_),
    .A2(_07792_),
    .B1(_07800_),
    .C1(_07797_),
    .X(_07838_));
 sky130_fd_sc_hd__nand2_1 _24749_ (.A(_07790_),
    .B(net738),
    .Y(_07839_));
 sky130_fd_sc_hd__o21ai_1 _24750_ (.A1(_07819_),
    .A2(_07838_),
    .B1(net739),
    .Y(_02284_));
 sky130_fd_sc_hd__clkbuf_8 _24751_ (.A(_09057_),
    .X(_07840_));
 sky130_fd_sc_hd__a211o_1 _24752_ (.A1(_02959_),
    .A2(_07792_),
    .B1(_07840_),
    .C1(_07801_),
    .X(_07841_));
 sky130_fd_sc_hd__nand2_1 _24753_ (.A(_07790_),
    .B(net878),
    .Y(_07842_));
 sky130_fd_sc_hd__o21ai_1 _24754_ (.A1(_07819_),
    .A2(_07841_),
    .B1(net879),
    .Y(_02285_));
 sky130_fd_sc_hd__a211o_1 _24755_ (.A1(_02963_),
    .A2(_07792_),
    .B1(_07840_),
    .C1(_07804_),
    .X(_07843_));
 sky130_fd_sc_hd__nand2_1 _24756_ (.A(_07790_),
    .B(net1430),
    .Y(_07844_));
 sky130_fd_sc_hd__o21ai_1 _24757_ (.A1(_07819_),
    .A2(_07843_),
    .B1(net1431),
    .Y(_02286_));
 sky130_fd_sc_hd__a211o_1 _24758_ (.A1(_02967_),
    .A2(_07792_),
    .B1(_07840_),
    .C1(_07807_),
    .X(_07845_));
 sky130_fd_sc_hd__nand2_1 _24759_ (.A(_07790_),
    .B(net834),
    .Y(_07846_));
 sky130_fd_sc_hd__o21ai_1 _24760_ (.A1(_07819_),
    .A2(_07845_),
    .B1(net835),
    .Y(_02287_));
 sky130_fd_sc_hd__a211o_1 _24761_ (.A1(_02971_),
    .A2(_07792_),
    .B1(_07840_),
    .C1(_07810_),
    .X(_07847_));
 sky130_fd_sc_hd__nand2_1 _24762_ (.A(_07790_),
    .B(net1306),
    .Y(_07848_));
 sky130_fd_sc_hd__o21ai_1 _24763_ (.A1(_07819_),
    .A2(_07847_),
    .B1(net1307),
    .Y(_02288_));
 sky130_fd_sc_hd__a211o_1 _24764_ (.A1(_02975_),
    .A2(_07792_),
    .B1(_07840_),
    .C1(_07813_),
    .X(_07849_));
 sky130_fd_sc_hd__nand2_1 _24765_ (.A(_07790_),
    .B(net746),
    .Y(_07850_));
 sky130_fd_sc_hd__o21ai_1 _24766_ (.A1(_07819_),
    .A2(_07849_),
    .B1(net747),
    .Y(_02289_));
 sky130_fd_sc_hd__a211o_1 _24767_ (.A1(_02979_),
    .A2(_07792_),
    .B1(_07840_),
    .C1(_07816_),
    .X(_07851_));
 sky130_fd_sc_hd__nand2_1 _24768_ (.A(_07790_),
    .B(net962),
    .Y(_07852_));
 sky130_fd_sc_hd__o21ai_1 _24769_ (.A1(_07819_),
    .A2(_07851_),
    .B1(net963),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _24770_ (.A(_03058_),
    .B(_09070_),
    .Y(_07853_));
 sky130_fd_sc_hd__inv_2 _24771_ (.A(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__o21ai_4 _24772_ (.A1(_06755_),
    .A2(_07854_),
    .B1(_12190_),
    .Y(_07855_));
 sky130_fd_sc_hd__mux2_1 _24773_ (.A0(_07699_),
    .A1(net2550),
    .S(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__clkbuf_1 _24774_ (.A(_07856_),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _24775_ (.A0(_07703_),
    .A1(net3788),
    .S(_07855_),
    .X(_07857_));
 sky130_fd_sc_hd__clkbuf_1 _24776_ (.A(_07857_),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _24777_ (.A0(_07705_),
    .A1(net3620),
    .S(_07855_),
    .X(_07858_));
 sky130_fd_sc_hd__clkbuf_1 _24778_ (.A(_07858_),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _24779_ (.A0(_07707_),
    .A1(net2100),
    .S(_07855_),
    .X(_07859_));
 sky130_fd_sc_hd__clkbuf_1 _24780_ (.A(_07859_),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _24781_ (.A0(_07709_),
    .A1(net3568),
    .S(_07855_),
    .X(_07860_));
 sky130_fd_sc_hd__clkbuf_1 _24782_ (.A(_07860_),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _24783_ (.A0(_07711_),
    .A1(net2179),
    .S(_07855_),
    .X(_07861_));
 sky130_fd_sc_hd__clkbuf_1 _24784_ (.A(_07861_),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _24785_ (.A0(_07713_),
    .A1(net3352),
    .S(_07855_),
    .X(_07862_));
 sky130_fd_sc_hd__clkbuf_1 _24786_ (.A(_07862_),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _24787_ (.A0(_07715_),
    .A1(net3091),
    .S(_07855_),
    .X(_07863_));
 sky130_fd_sc_hd__clkbuf_1 _24788_ (.A(_07863_),
    .X(_02298_));
 sky130_fd_sc_hd__buf_4 _24789_ (.A(_07855_),
    .X(_07864_));
 sky130_fd_sc_hd__buf_4 _24790_ (.A(_07854_),
    .X(_07865_));
 sky130_fd_sc_hd__buf_4 _24791_ (.A(_07854_),
    .X(_07866_));
 sky130_fd_sc_hd__nor2_1 _24792_ (.A(_12183_),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__a211o_1 _24793_ (.A1(_02851_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07867_),
    .X(_07868_));
 sky130_fd_sc_hd__buf_4 _24794_ (.A(_07855_),
    .X(_07869_));
 sky130_fd_sc_hd__nand2_1 _24795_ (.A(_07869_),
    .B(net1056),
    .Y(_07870_));
 sky130_fd_sc_hd__o21ai_1 _24796_ (.A1(_07864_),
    .A2(_07868_),
    .B1(net1057),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _24797_ (.A(_12196_),
    .B(_07866_),
    .Y(_07871_));
 sky130_fd_sc_hd__a211o_1 _24798_ (.A1(_02861_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07871_),
    .X(_07872_));
 sky130_fd_sc_hd__nand2_1 _24799_ (.A(_07869_),
    .B(net1404),
    .Y(_07873_));
 sky130_fd_sc_hd__o21ai_1 _24800_ (.A1(_07864_),
    .A2(_07872_),
    .B1(net1405),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _24801_ (.A(_12204_),
    .B(_07866_),
    .Y(_07874_));
 sky130_fd_sc_hd__a211o_1 _24802_ (.A1(_02868_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__nand2_1 _24803_ (.A(_07869_),
    .B(net1668),
    .Y(_07876_));
 sky130_fd_sc_hd__o21ai_1 _24804_ (.A1(_07864_),
    .A2(_07875_),
    .B1(net1669),
    .Y(_02301_));
 sky130_fd_sc_hd__nor2_1 _24805_ (.A(_12212_),
    .B(_07866_),
    .Y(_07877_));
 sky130_fd_sc_hd__a211o_1 _24806_ (.A1(_02875_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07877_),
    .X(_07878_));
 sky130_fd_sc_hd__nand2_1 _24807_ (.A(_07869_),
    .B(net1046),
    .Y(_07879_));
 sky130_fd_sc_hd__o21ai_1 _24808_ (.A1(_07864_),
    .A2(_07878_),
    .B1(net1047),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _24809_ (.A(_12220_),
    .B(_07866_),
    .Y(_07880_));
 sky130_fd_sc_hd__a211o_1 _24810_ (.A1(_02882_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__nand2_1 _24811_ (.A(_07869_),
    .B(net1220),
    .Y(_07882_));
 sky130_fd_sc_hd__o21ai_1 _24812_ (.A1(_07864_),
    .A2(_07881_),
    .B1(net1221),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _24813_ (.A(_12228_),
    .B(_07866_),
    .Y(_07883_));
 sky130_fd_sc_hd__a211o_1 _24814_ (.A1(_02889_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__nand2_1 _24815_ (.A(_07869_),
    .B(net926),
    .Y(_07885_));
 sky130_fd_sc_hd__o21ai_1 _24816_ (.A1(_07864_),
    .A2(_07884_),
    .B1(net927),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _24817_ (.A(_12236_),
    .B(_07866_),
    .Y(_07886_));
 sky130_fd_sc_hd__a211o_1 _24818_ (.A1(_02896_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07886_),
    .X(_07887_));
 sky130_fd_sc_hd__nand2_1 _24819_ (.A(_07869_),
    .B(net1182),
    .Y(_07888_));
 sky130_fd_sc_hd__o21ai_1 _24820_ (.A1(_07864_),
    .A2(_07887_),
    .B1(net1183),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _24821_ (.A(_12244_),
    .B(_07866_),
    .Y(_07889_));
 sky130_fd_sc_hd__a211o_1 _24822_ (.A1(_02903_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07889_),
    .X(_07890_));
 sky130_fd_sc_hd__nand2_1 _24823_ (.A(_07869_),
    .B(net1148),
    .Y(_07891_));
 sky130_fd_sc_hd__o21ai_1 _24824_ (.A1(_07864_),
    .A2(_07890_),
    .B1(net1149),
    .Y(_02306_));
 sky130_fd_sc_hd__buf_4 _24825_ (.A(_07855_),
    .X(_07892_));
 sky130_fd_sc_hd__a211o_1 _24826_ (.A1(_02911_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07867_),
    .X(_07893_));
 sky130_fd_sc_hd__nand2_1 _24827_ (.A(_07869_),
    .B(net1774),
    .Y(_07894_));
 sky130_fd_sc_hd__o21ai_1 _24828_ (.A1(_07892_),
    .A2(_07893_),
    .B1(net1775),
    .Y(_02307_));
 sky130_fd_sc_hd__a211o_1 _24829_ (.A1(_02916_),
    .A2(_07865_),
    .B1(_07840_),
    .C1(_07871_),
    .X(_07895_));
 sky130_fd_sc_hd__nand2_1 _24830_ (.A(_07869_),
    .B(net896),
    .Y(_07896_));
 sky130_fd_sc_hd__o21ai_1 _24831_ (.A1(_07892_),
    .A2(_07895_),
    .B1(net897),
    .Y(_02308_));
 sky130_fd_sc_hd__buf_4 _24832_ (.A(_09057_),
    .X(_07897_));
 sky130_fd_sc_hd__a211o_1 _24833_ (.A1(_02921_),
    .A2(_07865_),
    .B1(_07897_),
    .C1(_07874_),
    .X(_07898_));
 sky130_fd_sc_hd__nand2_1 _24834_ (.A(_07869_),
    .B(net958),
    .Y(_07899_));
 sky130_fd_sc_hd__o21ai_1 _24835_ (.A1(_07892_),
    .A2(_07898_),
    .B1(net959),
    .Y(_02309_));
 sky130_fd_sc_hd__a211o_1 _24836_ (.A1(_02927_),
    .A2(_07865_),
    .B1(_07897_),
    .C1(_07877_),
    .X(_07900_));
 sky130_fd_sc_hd__nand2_1 _24837_ (.A(_07869_),
    .B(net1578),
    .Y(_07901_));
 sky130_fd_sc_hd__o21ai_1 _24838_ (.A1(_07892_),
    .A2(_07900_),
    .B1(net1579),
    .Y(_02310_));
 sky130_fd_sc_hd__a211o_1 _24839_ (.A1(_02932_),
    .A2(_07865_),
    .B1(_07897_),
    .C1(_07880_),
    .X(_07902_));
 sky130_fd_sc_hd__nand2_1 _24840_ (.A(_07869_),
    .B(net1516),
    .Y(_07903_));
 sky130_fd_sc_hd__o21ai_1 _24841_ (.A1(_07892_),
    .A2(_07902_),
    .B1(net1517),
    .Y(_02311_));
 sky130_fd_sc_hd__a211o_1 _24842_ (.A1(_02937_),
    .A2(_07865_),
    .B1(_07897_),
    .C1(_07883_),
    .X(_07904_));
 sky130_fd_sc_hd__nand2_1 _24843_ (.A(_07869_),
    .B(net1262),
    .Y(_07905_));
 sky130_fd_sc_hd__o21ai_1 _24844_ (.A1(_07892_),
    .A2(_07904_),
    .B1(net1263),
    .Y(_02312_));
 sky130_fd_sc_hd__a211o_1 _24845_ (.A1(_02942_),
    .A2(_07865_),
    .B1(_07897_),
    .C1(_07886_),
    .X(_07906_));
 sky130_fd_sc_hd__nand2_1 _24846_ (.A(_07869_),
    .B(net1112),
    .Y(_07907_));
 sky130_fd_sc_hd__o21ai_1 _24847_ (.A1(_07892_),
    .A2(_07906_),
    .B1(net1113),
    .Y(_02313_));
 sky130_fd_sc_hd__a211o_1 _24848_ (.A1(_02947_),
    .A2(_07865_),
    .B1(_07897_),
    .C1(_07889_),
    .X(_07908_));
 sky130_fd_sc_hd__nand2_1 _24849_ (.A(_07869_),
    .B(net902),
    .Y(_07909_));
 sky130_fd_sc_hd__o21ai_1 _24850_ (.A1(_07892_),
    .A2(_07908_),
    .B1(net903),
    .Y(_02314_));
 sky130_fd_sc_hd__a211o_1 _24851_ (.A1(_02951_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07867_),
    .X(_07910_));
 sky130_fd_sc_hd__nand2_1 _24852_ (.A(_07864_),
    .B(net686),
    .Y(_07911_));
 sky130_fd_sc_hd__o21ai_1 _24853_ (.A1(_07892_),
    .A2(_07910_),
    .B1(net687),
    .Y(_02315_));
 sky130_fd_sc_hd__a211o_1 _24854_ (.A1(_02955_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07871_),
    .X(_07912_));
 sky130_fd_sc_hd__nand2_1 _24855_ (.A(_07864_),
    .B(net632),
    .Y(_07913_));
 sky130_fd_sc_hd__o21ai_1 _24856_ (.A1(_07892_),
    .A2(_07912_),
    .B1(net633),
    .Y(_02316_));
 sky130_fd_sc_hd__a211o_1 _24857_ (.A1(_02959_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07874_),
    .X(_07914_));
 sky130_fd_sc_hd__nand2_1 _24858_ (.A(_07864_),
    .B(net616),
    .Y(_07915_));
 sky130_fd_sc_hd__o21ai_1 _24859_ (.A1(_07892_),
    .A2(_07914_),
    .B1(net617),
    .Y(_02317_));
 sky130_fd_sc_hd__a211o_1 _24860_ (.A1(_02963_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07877_),
    .X(_07916_));
 sky130_fd_sc_hd__nand2_1 _24861_ (.A(_07864_),
    .B(net714),
    .Y(_07917_));
 sky130_fd_sc_hd__o21ai_1 _24862_ (.A1(_07892_),
    .A2(_07916_),
    .B1(net715),
    .Y(_02318_));
 sky130_fd_sc_hd__a211o_1 _24863_ (.A1(_02967_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07880_),
    .X(_07918_));
 sky130_fd_sc_hd__nand2_1 _24864_ (.A(_07864_),
    .B(net462),
    .Y(_07919_));
 sky130_fd_sc_hd__o21ai_1 _24865_ (.A1(_07892_),
    .A2(_07918_),
    .B1(net463),
    .Y(_02319_));
 sky130_fd_sc_hd__a211o_1 _24866_ (.A1(_02971_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07883_),
    .X(_07920_));
 sky130_fd_sc_hd__nand2_1 _24867_ (.A(_07864_),
    .B(net422),
    .Y(_07921_));
 sky130_fd_sc_hd__o21ai_1 _24868_ (.A1(_07892_),
    .A2(_07920_),
    .B1(net423),
    .Y(_02320_));
 sky130_fd_sc_hd__a211o_1 _24869_ (.A1(_02975_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07886_),
    .X(_07922_));
 sky130_fd_sc_hd__nand2_1 _24870_ (.A(_07864_),
    .B(net532),
    .Y(_07923_));
 sky130_fd_sc_hd__o21ai_1 _24871_ (.A1(_07892_),
    .A2(_07922_),
    .B1(net533),
    .Y(_02321_));
 sky130_fd_sc_hd__a211o_1 _24872_ (.A1(_02979_),
    .A2(_07866_),
    .B1(_07897_),
    .C1(_07889_),
    .X(_07924_));
 sky130_fd_sc_hd__nand2_1 _24873_ (.A(_07864_),
    .B(net488),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_1 _24874_ (.A1(_07892_),
    .A2(_07924_),
    .B1(net489),
    .Y(_02322_));
 sky130_fd_sc_hd__nor2_1 _24875_ (.A(_12313_),
    .B(_03133_),
    .Y(_07926_));
 sky130_fd_sc_hd__o21ai_4 _24876_ (.A1(_12289_),
    .A2(_07926_),
    .B1(_12190_),
    .Y(_07927_));
 sky130_fd_sc_hd__mux2_1 _24877_ (.A0(_07699_),
    .A1(net3425),
    .S(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__clkbuf_1 _24878_ (.A(_07928_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _24879_ (.A0(_07703_),
    .A1(net2680),
    .S(_07927_),
    .X(_07929_));
 sky130_fd_sc_hd__clkbuf_1 _24880_ (.A(_07929_),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _24881_ (.A0(_07705_),
    .A1(net2944),
    .S(_07927_),
    .X(_07930_));
 sky130_fd_sc_hd__clkbuf_1 _24882_ (.A(_07930_),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _24883_ (.A0(_07707_),
    .A1(net2340),
    .S(_07927_),
    .X(_07931_));
 sky130_fd_sc_hd__clkbuf_1 _24884_ (.A(_07931_),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _24885_ (.A0(_07709_),
    .A1(net2995),
    .S(_07927_),
    .X(_07932_));
 sky130_fd_sc_hd__clkbuf_1 _24886_ (.A(_07932_),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _24887_ (.A0(_07711_),
    .A1(net3547),
    .S(_07927_),
    .X(_07933_));
 sky130_fd_sc_hd__clkbuf_1 _24888_ (.A(_07933_),
    .X(_02328_));
 sky130_fd_sc_hd__mux2_1 _24889_ (.A0(_07713_),
    .A1(net3665),
    .S(_07927_),
    .X(_07934_));
 sky130_fd_sc_hd__clkbuf_1 _24890_ (.A(_07934_),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _24891_ (.A0(_07715_),
    .A1(net3518),
    .S(_07927_),
    .X(_07935_));
 sky130_fd_sc_hd__clkbuf_1 _24892_ (.A(_07935_),
    .X(_02330_));
 sky130_fd_sc_hd__buf_4 _24893_ (.A(_07927_),
    .X(_07936_));
 sky130_fd_sc_hd__buf_4 _24894_ (.A(_07926_),
    .X(_07937_));
 sky130_fd_sc_hd__buf_4 _24895_ (.A(_07926_),
    .X(_07938_));
 sky130_fd_sc_hd__nor2_1 _24896_ (.A(_12183_),
    .B(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__a211o_1 _24897_ (.A1(_02851_),
    .A2(_07937_),
    .B1(_07897_),
    .C1(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__buf_4 _24898_ (.A(_07927_),
    .X(_07941_));
 sky130_fd_sc_hd__nand2_1 _24899_ (.A(_07941_),
    .B(net1298),
    .Y(_07942_));
 sky130_fd_sc_hd__o21ai_1 _24900_ (.A1(_07936_),
    .A2(_07940_),
    .B1(net1299),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _24901_ (.A(_12196_),
    .B(_07938_),
    .Y(_07943_));
 sky130_fd_sc_hd__a211o_1 _24902_ (.A1(_02861_),
    .A2(_07937_),
    .B1(_07897_),
    .C1(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__nand2_1 _24903_ (.A(_07941_),
    .B(net1899),
    .Y(_07945_));
 sky130_fd_sc_hd__o21ai_1 _24904_ (.A1(_07936_),
    .A2(_07944_),
    .B1(net1900),
    .Y(_02332_));
 sky130_fd_sc_hd__buf_4 _24905_ (.A(_09057_),
    .X(_07946_));
 sky130_fd_sc_hd__nor2_1 _24906_ (.A(_12204_),
    .B(_07938_),
    .Y(_07947_));
 sky130_fd_sc_hd__a211o_1 _24907_ (.A1(_02868_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__nand2_1 _24908_ (.A(_07941_),
    .B(net1532),
    .Y(_07949_));
 sky130_fd_sc_hd__o21ai_1 _24909_ (.A1(_07936_),
    .A2(_07948_),
    .B1(net1533),
    .Y(_02333_));
 sky130_fd_sc_hd__nor2_1 _24910_ (.A(_12212_),
    .B(_07938_),
    .Y(_07950_));
 sky130_fd_sc_hd__a211o_1 _24911_ (.A1(_02875_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07950_),
    .X(_07951_));
 sky130_fd_sc_hd__nand2_1 _24912_ (.A(_07941_),
    .B(net1612),
    .Y(_07952_));
 sky130_fd_sc_hd__o21ai_1 _24913_ (.A1(_07936_),
    .A2(_07951_),
    .B1(net1613),
    .Y(_02334_));
 sky130_fd_sc_hd__nor2_1 _24914_ (.A(_12220_),
    .B(_07938_),
    .Y(_07953_));
 sky130_fd_sc_hd__a211o_1 _24915_ (.A1(_02882_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__nand2_1 _24916_ (.A(_07941_),
    .B(net1384),
    .Y(_07955_));
 sky130_fd_sc_hd__o21ai_1 _24917_ (.A1(_07936_),
    .A2(_07954_),
    .B1(net1385),
    .Y(_02335_));
 sky130_fd_sc_hd__nor2_1 _24918_ (.A(_12228_),
    .B(_07938_),
    .Y(_07956_));
 sky130_fd_sc_hd__a211o_1 _24919_ (.A1(_02889_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07956_),
    .X(_07957_));
 sky130_fd_sc_hd__nand2_1 _24920_ (.A(_07941_),
    .B(net1614),
    .Y(_07958_));
 sky130_fd_sc_hd__o21ai_1 _24921_ (.A1(_07936_),
    .A2(_07957_),
    .B1(net1615),
    .Y(_02336_));
 sky130_fd_sc_hd__nor2_1 _24922_ (.A(_12236_),
    .B(_07938_),
    .Y(_07959_));
 sky130_fd_sc_hd__a211o_1 _24923_ (.A1(_02896_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__nand2_1 _24924_ (.A(_07941_),
    .B(net970),
    .Y(_07961_));
 sky130_fd_sc_hd__o21ai_1 _24925_ (.A1(_07936_),
    .A2(_07960_),
    .B1(net971),
    .Y(_02337_));
 sky130_fd_sc_hd__nor2_1 _24926_ (.A(_12244_),
    .B(_07938_),
    .Y(_07962_));
 sky130_fd_sc_hd__a211o_1 _24927_ (.A1(_02903_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__nand2_1 _24928_ (.A(_07941_),
    .B(net1656),
    .Y(_07964_));
 sky130_fd_sc_hd__o21ai_1 _24929_ (.A1(_07936_),
    .A2(_07963_),
    .B1(net1657),
    .Y(_02338_));
 sky130_fd_sc_hd__buf_4 _24930_ (.A(_07927_),
    .X(_07965_));
 sky130_fd_sc_hd__a211o_1 _24931_ (.A1(_02911_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07939_),
    .X(_07966_));
 sky130_fd_sc_hd__nand2_1 _24932_ (.A(_07941_),
    .B(net1420),
    .Y(_07967_));
 sky130_fd_sc_hd__o21ai_1 _24933_ (.A1(_07965_),
    .A2(_07966_),
    .B1(net1421),
    .Y(_02339_));
 sky130_fd_sc_hd__a211o_1 _24934_ (.A1(_02916_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07943_),
    .X(_07968_));
 sky130_fd_sc_hd__nand2_1 _24935_ (.A(_07941_),
    .B(net1844),
    .Y(_07969_));
 sky130_fd_sc_hd__o21ai_1 _24936_ (.A1(_07965_),
    .A2(_07968_),
    .B1(net1845),
    .Y(_02340_));
 sky130_fd_sc_hd__a211o_1 _24937_ (.A1(_02921_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07947_),
    .X(_07970_));
 sky130_fd_sc_hd__nand2_1 _24938_ (.A(_07941_),
    .B(net1048),
    .Y(_07971_));
 sky130_fd_sc_hd__o21ai_1 _24939_ (.A1(_07965_),
    .A2(_07970_),
    .B1(net1049),
    .Y(_02341_));
 sky130_fd_sc_hd__a211o_1 _24940_ (.A1(_02927_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07950_),
    .X(_07972_));
 sky130_fd_sc_hd__nand2_1 _24941_ (.A(_07941_),
    .B(net1696),
    .Y(_07973_));
 sky130_fd_sc_hd__o21ai_1 _24942_ (.A1(_07965_),
    .A2(_07972_),
    .B1(net1697),
    .Y(_02342_));
 sky130_fd_sc_hd__a211o_1 _24943_ (.A1(_02932_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07953_),
    .X(_07974_));
 sky130_fd_sc_hd__nand2_1 _24944_ (.A(_07941_),
    .B(net1514),
    .Y(_07975_));
 sky130_fd_sc_hd__o21ai_1 _24945_ (.A1(_07965_),
    .A2(_07974_),
    .B1(net1515),
    .Y(_02343_));
 sky130_fd_sc_hd__a211o_1 _24946_ (.A1(_02937_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07956_),
    .X(_07976_));
 sky130_fd_sc_hd__nand2_1 _24947_ (.A(_07941_),
    .B(net1576),
    .Y(_07977_));
 sky130_fd_sc_hd__o21ai_1 _24948_ (.A1(_07965_),
    .A2(_07976_),
    .B1(net1577),
    .Y(_02344_));
 sky130_fd_sc_hd__a211o_1 _24949_ (.A1(_02942_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07959_),
    .X(_07978_));
 sky130_fd_sc_hd__nand2_1 _24950_ (.A(_07941_),
    .B(net1218),
    .Y(_07979_));
 sky130_fd_sc_hd__o21ai_1 _24951_ (.A1(_07965_),
    .A2(_07978_),
    .B1(net1219),
    .Y(_02345_));
 sky130_fd_sc_hd__a211o_1 _24952_ (.A1(_02947_),
    .A2(_07937_),
    .B1(_07946_),
    .C1(_07962_),
    .X(_07980_));
 sky130_fd_sc_hd__nand2_1 _24953_ (.A(_07941_),
    .B(net1536),
    .Y(_07981_));
 sky130_fd_sc_hd__o21ai_1 _24954_ (.A1(_07965_),
    .A2(_07980_),
    .B1(net1537),
    .Y(_02346_));
 sky130_fd_sc_hd__a211o_1 _24955_ (.A1(_02951_),
    .A2(_07938_),
    .B1(_07946_),
    .C1(_07939_),
    .X(_07982_));
 sky130_fd_sc_hd__nand2_1 _24956_ (.A(_07936_),
    .B(net1362),
    .Y(_07983_));
 sky130_fd_sc_hd__o21ai_1 _24957_ (.A1(_07965_),
    .A2(_07982_),
    .B1(net1363),
    .Y(_02347_));
 sky130_fd_sc_hd__a211o_1 _24958_ (.A1(_02955_),
    .A2(_07938_),
    .B1(_07946_),
    .C1(_07943_),
    .X(_07984_));
 sky130_fd_sc_hd__nand2_1 _24959_ (.A(_07936_),
    .B(net952),
    .Y(_07985_));
 sky130_fd_sc_hd__o21ai_1 _24960_ (.A1(_07965_),
    .A2(_07984_),
    .B1(net953),
    .Y(_02348_));
 sky130_fd_sc_hd__a211o_1 _24961_ (.A1(_02959_),
    .A2(_07938_),
    .B1(_12851_),
    .C1(_07947_),
    .X(_07986_));
 sky130_fd_sc_hd__nand2_1 _24962_ (.A(_07936_),
    .B(net838),
    .Y(_07987_));
 sky130_fd_sc_hd__o21ai_1 _24963_ (.A1(_07965_),
    .A2(_07986_),
    .B1(net839),
    .Y(_02349_));
 sky130_fd_sc_hd__a211o_1 _24964_ (.A1(_02963_),
    .A2(_07938_),
    .B1(_12851_),
    .C1(_07950_),
    .X(_07988_));
 sky130_fd_sc_hd__nand2_1 _24965_ (.A(_07936_),
    .B(net676),
    .Y(_07989_));
 sky130_fd_sc_hd__o21ai_1 _24966_ (.A1(_07965_),
    .A2(_07988_),
    .B1(net677),
    .Y(_02350_));
 sky130_fd_sc_hd__a211o_1 _24967_ (.A1(_02967_),
    .A2(_07938_),
    .B1(_12851_),
    .C1(_07953_),
    .X(_07990_));
 sky130_fd_sc_hd__nand2_1 _24968_ (.A(_07936_),
    .B(net716),
    .Y(_07991_));
 sky130_fd_sc_hd__o21ai_1 _24969_ (.A1(_07965_),
    .A2(_07990_),
    .B1(net717),
    .Y(_02351_));
 sky130_fd_sc_hd__a211o_1 _24970_ (.A1(_02971_),
    .A2(_07938_),
    .B1(_12851_),
    .C1(_07956_),
    .X(_07992_));
 sky130_fd_sc_hd__nand2_1 _24971_ (.A(_07936_),
    .B(net828),
    .Y(_07993_));
 sky130_fd_sc_hd__o21ai_1 _24972_ (.A1(_07965_),
    .A2(_07992_),
    .B1(net829),
    .Y(_02352_));
 sky130_fd_sc_hd__a211o_1 _24973_ (.A1(_02975_),
    .A2(_07938_),
    .B1(_12851_),
    .C1(_07959_),
    .X(_07994_));
 sky130_fd_sc_hd__nand2_1 _24974_ (.A(_07936_),
    .B(net598),
    .Y(_07995_));
 sky130_fd_sc_hd__o21ai_1 _24975_ (.A1(_07965_),
    .A2(_07994_),
    .B1(net599),
    .Y(_02353_));
 sky130_fd_sc_hd__a211o_1 _24976_ (.A1(_02979_),
    .A2(_07938_),
    .B1(_12851_),
    .C1(_07962_),
    .X(_07996_));
 sky130_fd_sc_hd__nand2_1 _24977_ (.A(_07936_),
    .B(net886),
    .Y(_07997_));
 sky130_fd_sc_hd__o21ai_1 _24978_ (.A1(_07965_),
    .A2(_07996_),
    .B1(net887),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _24979_ (.A(_03210_),
    .B(_12177_),
    .Y(_07998_));
 sky130_fd_sc_hd__a21bo_1 _24980_ (.A1(_07998_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_07999_));
 sky130_fd_sc_hd__clkbuf_8 _24981_ (.A(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__mux2_1 _24982_ (.A0(_07699_),
    .A1(net2885),
    .S(_08000_),
    .X(_08001_));
 sky130_fd_sc_hd__clkbuf_1 _24983_ (.A(_08001_),
    .X(_02355_));
 sky130_fd_sc_hd__mux2_1 _24984_ (.A0(_07703_),
    .A1(net2764),
    .S(_08000_),
    .X(_08002_));
 sky130_fd_sc_hd__clkbuf_1 _24985_ (.A(_08002_),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _24986_ (.A0(_07705_),
    .A1(net3174),
    .S(_08000_),
    .X(_08003_));
 sky130_fd_sc_hd__clkbuf_1 _24987_ (.A(_08003_),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _24988_ (.A0(_07707_),
    .A1(net3541),
    .S(_08000_),
    .X(_08004_));
 sky130_fd_sc_hd__clkbuf_1 _24989_ (.A(_08004_),
    .X(_02358_));
 sky130_fd_sc_hd__mux2_1 _24990_ (.A0(_07709_),
    .A1(net3292),
    .S(_08000_),
    .X(_08005_));
 sky130_fd_sc_hd__clkbuf_1 _24991_ (.A(_08005_),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _24992_ (.A0(_07711_),
    .A1(net2853),
    .S(_08000_),
    .X(_08006_));
 sky130_fd_sc_hd__clkbuf_1 _24993_ (.A(_08006_),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _24994_ (.A0(_07713_),
    .A1(net2613),
    .S(_08000_),
    .X(_08007_));
 sky130_fd_sc_hd__clkbuf_1 _24995_ (.A(_08007_),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _24996_ (.A0(_07715_),
    .A1(net3483),
    .S(_08000_),
    .X(_08008_));
 sky130_fd_sc_hd__clkbuf_1 _24997_ (.A(_08008_),
    .X(_02362_));
 sky130_fd_sc_hd__buf_4 _24998_ (.A(_07998_),
    .X(_08009_));
 sky130_fd_sc_hd__buf_4 _24999_ (.A(_06885_),
    .X(_08010_));
 sky130_fd_sc_hd__buf_4 _25000_ (.A(_07998_),
    .X(_08011_));
 sky130_fd_sc_hd__nand2_1 _25001_ (.A(_08011_),
    .B(_12184_),
    .Y(_08012_));
 sky130_fd_sc_hd__o211a_1 _25002_ (.A1(_02850_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__mux2_1 _25003_ (.A0(_08013_),
    .A1(net3279),
    .S(_08000_),
    .X(_08014_));
 sky130_fd_sc_hd__clkbuf_1 _25004_ (.A(_08014_),
    .X(_02363_));
 sky130_fd_sc_hd__nand2_1 _25005_ (.A(_08011_),
    .B(_12197_),
    .Y(_08015_));
 sky130_fd_sc_hd__o211a_1 _25006_ (.A1(_02860_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__mux2_1 _25007_ (.A0(_08016_),
    .A1(net2957),
    .S(_08000_),
    .X(_08017_));
 sky130_fd_sc_hd__clkbuf_1 _25008_ (.A(_08017_),
    .X(_02364_));
 sky130_fd_sc_hd__nand2_1 _25009_ (.A(_08011_),
    .B(_12205_),
    .Y(_08018_));
 sky130_fd_sc_hd__o211a_1 _25010_ (.A1(_02867_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08018_),
    .X(_08019_));
 sky130_fd_sc_hd__mux2_1 _25011_ (.A0(_08019_),
    .A1(net2491),
    .S(_08000_),
    .X(_08020_));
 sky130_fd_sc_hd__clkbuf_1 _25012_ (.A(_08020_),
    .X(_02365_));
 sky130_fd_sc_hd__nand2_1 _25013_ (.A(_08011_),
    .B(_12213_),
    .Y(_08021_));
 sky130_fd_sc_hd__o211a_1 _25014_ (.A1(_02874_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08021_),
    .X(_08022_));
 sky130_fd_sc_hd__mux2_1 _25015_ (.A0(_08022_),
    .A1(net3136),
    .S(_08000_),
    .X(_08023_));
 sky130_fd_sc_hd__clkbuf_1 _25016_ (.A(_08023_),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_1 _25017_ (.A(_08011_),
    .B(_12221_),
    .Y(_08024_));
 sky130_fd_sc_hd__o211a_1 _25018_ (.A1(_02881_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__mux2_1 _25019_ (.A0(_08025_),
    .A1(net2692),
    .S(_08000_),
    .X(_08026_));
 sky130_fd_sc_hd__clkbuf_1 _25020_ (.A(_08026_),
    .X(_02367_));
 sky130_fd_sc_hd__nand2_1 _25021_ (.A(_08011_),
    .B(_12229_),
    .Y(_08027_));
 sky130_fd_sc_hd__o211a_1 _25022_ (.A1(_02888_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__mux2_1 _25023_ (.A0(_08028_),
    .A1(net2264),
    .S(_08000_),
    .X(_08029_));
 sky130_fd_sc_hd__clkbuf_1 _25024_ (.A(_08029_),
    .X(_02368_));
 sky130_fd_sc_hd__nand2_1 _25025_ (.A(_08011_),
    .B(_12237_),
    .Y(_08030_));
 sky130_fd_sc_hd__o211a_1 _25026_ (.A1(_02895_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__mux2_1 _25027_ (.A0(_08031_),
    .A1(net2430),
    .S(_08000_),
    .X(_08032_));
 sky130_fd_sc_hd__clkbuf_1 _25028_ (.A(_08032_),
    .X(_02369_));
 sky130_fd_sc_hd__nand2_1 _25029_ (.A(_08011_),
    .B(_12245_),
    .Y(_08033_));
 sky130_fd_sc_hd__o211a_1 _25030_ (.A1(_02902_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__mux2_1 _25031_ (.A0(_08034_),
    .A1(net2526),
    .S(_08000_),
    .X(_08035_));
 sky130_fd_sc_hd__clkbuf_1 _25032_ (.A(_08035_),
    .X(_02370_));
 sky130_fd_sc_hd__o211a_1 _25033_ (.A1(_02910_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08012_),
    .X(_08036_));
 sky130_fd_sc_hd__clkbuf_8 _25034_ (.A(_07999_),
    .X(_08037_));
 sky130_fd_sc_hd__mux2_1 _25035_ (.A0(_08036_),
    .A1(net2689),
    .S(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__clkbuf_1 _25036_ (.A(_08038_),
    .X(_02371_));
 sky130_fd_sc_hd__o211a_1 _25037_ (.A1(_02915_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08015_),
    .X(_08039_));
 sky130_fd_sc_hd__mux2_1 _25038_ (.A0(_08039_),
    .A1(net3485),
    .S(_08037_),
    .X(_08040_));
 sky130_fd_sc_hd__clkbuf_1 _25039_ (.A(_08040_),
    .X(_02372_));
 sky130_fd_sc_hd__o211a_1 _25040_ (.A1(_02920_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08018_),
    .X(_08041_));
 sky130_fd_sc_hd__mux2_1 _25041_ (.A0(_08041_),
    .A1(net3064),
    .S(_08037_),
    .X(_08042_));
 sky130_fd_sc_hd__clkbuf_1 _25042_ (.A(_08042_),
    .X(_02373_));
 sky130_fd_sc_hd__o211a_1 _25043_ (.A1(_02926_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08021_),
    .X(_08043_));
 sky130_fd_sc_hd__mux2_1 _25044_ (.A0(_08043_),
    .A1(net3561),
    .S(_08037_),
    .X(_08044_));
 sky130_fd_sc_hd__clkbuf_1 _25045_ (.A(_08044_),
    .X(_02374_));
 sky130_fd_sc_hd__o211a_1 _25046_ (.A1(_02931_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08024_),
    .X(_08045_));
 sky130_fd_sc_hd__mux2_1 _25047_ (.A0(_08045_),
    .A1(net3435),
    .S(_08037_),
    .X(_08046_));
 sky130_fd_sc_hd__clkbuf_1 _25048_ (.A(_08046_),
    .X(_02375_));
 sky130_fd_sc_hd__o211a_1 _25049_ (.A1(_02936_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08027_),
    .X(_08047_));
 sky130_fd_sc_hd__mux2_1 _25050_ (.A0(_08047_),
    .A1(net2722),
    .S(_08037_),
    .X(_08048_));
 sky130_fd_sc_hd__clkbuf_1 _25051_ (.A(_08048_),
    .X(_02376_));
 sky130_fd_sc_hd__o211a_1 _25052_ (.A1(_02941_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08030_),
    .X(_08049_));
 sky130_fd_sc_hd__mux2_1 _25053_ (.A0(_08049_),
    .A1(net2630),
    .S(_08037_),
    .X(_08050_));
 sky130_fd_sc_hd__clkbuf_1 _25054_ (.A(_08050_),
    .X(_02377_));
 sky130_fd_sc_hd__o211a_1 _25055_ (.A1(_02946_),
    .A2(_08009_),
    .B1(_08010_),
    .C1(_08033_),
    .X(_08051_));
 sky130_fd_sc_hd__mux2_1 _25056_ (.A0(_08051_),
    .A1(net2312),
    .S(_08037_),
    .X(_08052_));
 sky130_fd_sc_hd__clkbuf_1 _25057_ (.A(_08052_),
    .X(_02378_));
 sky130_fd_sc_hd__buf_4 _25058_ (.A(_06885_),
    .X(_08053_));
 sky130_fd_sc_hd__o211a_1 _25059_ (.A1(_12169_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08012_),
    .X(_08054_));
 sky130_fd_sc_hd__mux2_1 _25060_ (.A0(_08054_),
    .A1(net2817),
    .S(_08037_),
    .X(_08055_));
 sky130_fd_sc_hd__clkbuf_1 _25061_ (.A(_08055_),
    .X(_02379_));
 sky130_fd_sc_hd__o211a_1 _25062_ (.A1(_12194_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08015_),
    .X(_08056_));
 sky130_fd_sc_hd__mux2_1 _25063_ (.A0(_08056_),
    .A1(net3496),
    .S(_08037_),
    .X(_08057_));
 sky130_fd_sc_hd__clkbuf_1 _25064_ (.A(_08057_),
    .X(_02380_));
 sky130_fd_sc_hd__o211a_1 _25065_ (.A1(_12202_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08018_),
    .X(_08058_));
 sky130_fd_sc_hd__mux2_1 _25066_ (.A0(_08058_),
    .A1(net2444),
    .S(_08037_),
    .X(_08059_));
 sky130_fd_sc_hd__clkbuf_1 _25067_ (.A(_08059_),
    .X(_02381_));
 sky130_fd_sc_hd__o211a_1 _25068_ (.A1(_12210_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08021_),
    .X(_08060_));
 sky130_fd_sc_hd__mux2_1 _25069_ (.A0(_08060_),
    .A1(net2315),
    .S(_08037_),
    .X(_08061_));
 sky130_fd_sc_hd__clkbuf_1 _25070_ (.A(_08061_),
    .X(_02382_));
 sky130_fd_sc_hd__o211a_1 _25071_ (.A1(_12218_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08024_),
    .X(_08062_));
 sky130_fd_sc_hd__mux2_1 _25072_ (.A0(_08062_),
    .A1(net2349),
    .S(_08037_),
    .X(_08063_));
 sky130_fd_sc_hd__clkbuf_1 _25073_ (.A(_08063_),
    .X(_02383_));
 sky130_fd_sc_hd__o211a_1 _25074_ (.A1(_12226_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08027_),
    .X(_08064_));
 sky130_fd_sc_hd__mux2_1 _25075_ (.A0(_08064_),
    .A1(net2823),
    .S(_08037_),
    .X(_08065_));
 sky130_fd_sc_hd__clkbuf_1 _25076_ (.A(_08065_),
    .X(_02384_));
 sky130_fd_sc_hd__o211a_1 _25077_ (.A1(_12234_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08030_),
    .X(_08066_));
 sky130_fd_sc_hd__mux2_1 _25078_ (.A0(_08066_),
    .A1(net2850),
    .S(_08037_),
    .X(_08067_));
 sky130_fd_sc_hd__clkbuf_1 _25079_ (.A(_08067_),
    .X(_02385_));
 sky130_fd_sc_hd__o211a_1 _25080_ (.A1(_12242_),
    .A2(_08011_),
    .B1(_08053_),
    .C1(_08033_),
    .X(_08068_));
 sky130_fd_sc_hd__mux2_1 _25081_ (.A0(_08068_),
    .A1(net2342),
    .S(_08037_),
    .X(_08069_));
 sky130_fd_sc_hd__clkbuf_1 _25082_ (.A(_08069_),
    .X(_02386_));
 sky130_fd_sc_hd__nand2_1 _25083_ (.A(_03298_),
    .B(_12177_),
    .Y(_08070_));
 sky130_fd_sc_hd__a21bo_1 _25084_ (.A1(_08070_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_08071_));
 sky130_fd_sc_hd__clkbuf_8 _25085_ (.A(_08071_),
    .X(_08072_));
 sky130_fd_sc_hd__mux2_1 _25086_ (.A0(_07699_),
    .A1(net2511),
    .S(_08072_),
    .X(_08073_));
 sky130_fd_sc_hd__clkbuf_1 _25087_ (.A(_08073_),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _25088_ (.A0(_07703_),
    .A1(net2591),
    .S(_08072_),
    .X(_08074_));
 sky130_fd_sc_hd__clkbuf_1 _25089_ (.A(_08074_),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _25090_ (.A0(_07705_),
    .A1(net3197),
    .S(_08072_),
    .X(_08075_));
 sky130_fd_sc_hd__clkbuf_1 _25091_ (.A(_08075_),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _25092_ (.A0(_07707_),
    .A1(net3387),
    .S(_08072_),
    .X(_08076_));
 sky130_fd_sc_hd__clkbuf_1 _25093_ (.A(_08076_),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _25094_ (.A0(_07709_),
    .A1(net2299),
    .S(_08072_),
    .X(_08077_));
 sky130_fd_sc_hd__clkbuf_1 _25095_ (.A(_08077_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _25096_ (.A0(_07711_),
    .A1(net2674),
    .S(_08072_),
    .X(_08078_));
 sky130_fd_sc_hd__clkbuf_1 _25097_ (.A(_08078_),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _25098_ (.A0(_07713_),
    .A1(net2502),
    .S(_08072_),
    .X(_08079_));
 sky130_fd_sc_hd__clkbuf_1 _25099_ (.A(_08079_),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _25100_ (.A0(_07715_),
    .A1(net3042),
    .S(_08072_),
    .X(_08080_));
 sky130_fd_sc_hd__clkbuf_1 _25101_ (.A(_08080_),
    .X(_02394_));
 sky130_fd_sc_hd__buf_4 _25102_ (.A(_08070_),
    .X(_08081_));
 sky130_fd_sc_hd__buf_4 _25103_ (.A(_08070_),
    .X(_08082_));
 sky130_fd_sc_hd__nand2_1 _25104_ (.A(_08082_),
    .B(_12184_),
    .Y(_08083_));
 sky130_fd_sc_hd__o211a_1 _25105_ (.A1(_02850_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__mux2_1 _25106_ (.A0(_08084_),
    .A1(net3413),
    .S(_08072_),
    .X(_08085_));
 sky130_fd_sc_hd__clkbuf_1 _25107_ (.A(_08085_),
    .X(_02395_));
 sky130_fd_sc_hd__nand2_1 _25108_ (.A(_08082_),
    .B(_12197_),
    .Y(_08086_));
 sky130_fd_sc_hd__o211a_1 _25109_ (.A1(_02860_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08086_),
    .X(_08087_));
 sky130_fd_sc_hd__mux2_1 _25110_ (.A0(_08087_),
    .A1(net3474),
    .S(_08072_),
    .X(_08088_));
 sky130_fd_sc_hd__clkbuf_1 _25111_ (.A(_08088_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_1 _25112_ (.A(_08082_),
    .B(_12205_),
    .Y(_08089_));
 sky130_fd_sc_hd__o211a_1 _25113_ (.A1(_02867_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__mux2_1 _25114_ (.A0(_08090_),
    .A1(net2605),
    .S(_08072_),
    .X(_08091_));
 sky130_fd_sc_hd__clkbuf_1 _25115_ (.A(_08091_),
    .X(_02397_));
 sky130_fd_sc_hd__nand2_1 _25116_ (.A(_08082_),
    .B(_12213_),
    .Y(_08092_));
 sky130_fd_sc_hd__o211a_1 _25117_ (.A1(_02874_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__mux2_1 _25118_ (.A0(_08093_),
    .A1(net2481),
    .S(_08072_),
    .X(_08094_));
 sky130_fd_sc_hd__clkbuf_1 _25119_ (.A(_08094_),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_1 _25120_ (.A(_08082_),
    .B(_12221_),
    .Y(_08095_));
 sky130_fd_sc_hd__o211a_1 _25121_ (.A1(_02881_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__mux2_1 _25122_ (.A0(_08096_),
    .A1(net2787),
    .S(_08072_),
    .X(_08097_));
 sky130_fd_sc_hd__clkbuf_1 _25123_ (.A(_08097_),
    .X(_02399_));
 sky130_fd_sc_hd__nand2_1 _25124_ (.A(_08082_),
    .B(_12229_),
    .Y(_08098_));
 sky130_fd_sc_hd__o211a_1 _25125_ (.A1(_02888_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08098_),
    .X(_08099_));
 sky130_fd_sc_hd__mux2_1 _25126_ (.A0(_08099_),
    .A1(net3123),
    .S(_08072_),
    .X(_08100_));
 sky130_fd_sc_hd__clkbuf_1 _25127_ (.A(_08100_),
    .X(_02400_));
 sky130_fd_sc_hd__nand2_1 _25128_ (.A(_08082_),
    .B(_12237_),
    .Y(_08101_));
 sky130_fd_sc_hd__o211a_1 _25129_ (.A1(_02895_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08101_),
    .X(_08102_));
 sky130_fd_sc_hd__mux2_1 _25130_ (.A0(_08102_),
    .A1(net3529),
    .S(_08072_),
    .X(_08103_));
 sky130_fd_sc_hd__clkbuf_1 _25131_ (.A(_08103_),
    .X(_02401_));
 sky130_fd_sc_hd__nand2_1 _25132_ (.A(_08082_),
    .B(_12245_),
    .Y(_08104_));
 sky130_fd_sc_hd__o211a_1 _25133_ (.A1(_02902_),
    .A2(_08081_),
    .B1(_08053_),
    .C1(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__mux2_1 _25134_ (.A0(_08105_),
    .A1(net3427),
    .S(_08072_),
    .X(_08106_));
 sky130_fd_sc_hd__clkbuf_1 _25135_ (.A(_08106_),
    .X(_02402_));
 sky130_fd_sc_hd__buf_4 _25136_ (.A(_06885_),
    .X(_08107_));
 sky130_fd_sc_hd__o211a_1 _25137_ (.A1(_02910_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08083_),
    .X(_08108_));
 sky130_fd_sc_hd__clkbuf_8 _25138_ (.A(_08071_),
    .X(_08109_));
 sky130_fd_sc_hd__mux2_1 _25139_ (.A0(_08108_),
    .A1(net2159),
    .S(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__clkbuf_1 _25140_ (.A(_08110_),
    .X(_02403_));
 sky130_fd_sc_hd__o211a_1 _25141_ (.A1(_02915_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08086_),
    .X(_08111_));
 sky130_fd_sc_hd__mux2_1 _25142_ (.A0(_08111_),
    .A1(net2964),
    .S(_08109_),
    .X(_08112_));
 sky130_fd_sc_hd__clkbuf_1 _25143_ (.A(_08112_),
    .X(_02404_));
 sky130_fd_sc_hd__o211a_1 _25144_ (.A1(_02920_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08089_),
    .X(_08113_));
 sky130_fd_sc_hd__mux2_1 _25145_ (.A0(_08113_),
    .A1(net2503),
    .S(_08109_),
    .X(_08114_));
 sky130_fd_sc_hd__clkbuf_1 _25146_ (.A(_08114_),
    .X(_02405_));
 sky130_fd_sc_hd__o211a_1 _25147_ (.A1(_02926_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08092_),
    .X(_08115_));
 sky130_fd_sc_hd__mux2_1 _25148_ (.A0(_08115_),
    .A1(net3085),
    .S(_08109_),
    .X(_08116_));
 sky130_fd_sc_hd__clkbuf_1 _25149_ (.A(_08116_),
    .X(_02406_));
 sky130_fd_sc_hd__o211a_1 _25150_ (.A1(_02931_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08095_),
    .X(_08117_));
 sky130_fd_sc_hd__mux2_1 _25151_ (.A0(_08117_),
    .A1(net2509),
    .S(_08109_),
    .X(_08118_));
 sky130_fd_sc_hd__clkbuf_1 _25152_ (.A(_08118_),
    .X(_02407_));
 sky130_fd_sc_hd__o211a_1 _25153_ (.A1(_02936_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08098_),
    .X(_08119_));
 sky130_fd_sc_hd__mux2_1 _25154_ (.A0(_08119_),
    .A1(net2585),
    .S(_08109_),
    .X(_08120_));
 sky130_fd_sc_hd__clkbuf_1 _25155_ (.A(_08120_),
    .X(_02408_));
 sky130_fd_sc_hd__o211a_1 _25156_ (.A1(_02941_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08101_),
    .X(_08121_));
 sky130_fd_sc_hd__mux2_1 _25157_ (.A0(_08121_),
    .A1(net3092),
    .S(_08109_),
    .X(_08122_));
 sky130_fd_sc_hd__clkbuf_1 _25158_ (.A(_08122_),
    .X(_02409_));
 sky130_fd_sc_hd__o211a_1 _25159_ (.A1(_02946_),
    .A2(_08081_),
    .B1(_08107_),
    .C1(_08104_),
    .X(_08123_));
 sky130_fd_sc_hd__mux2_1 _25160_ (.A0(_08123_),
    .A1(net2380),
    .S(_08109_),
    .X(_08124_));
 sky130_fd_sc_hd__clkbuf_1 _25161_ (.A(_08124_),
    .X(_02410_));
 sky130_fd_sc_hd__o211a_1 _25162_ (.A1(_12169_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08083_),
    .X(_08125_));
 sky130_fd_sc_hd__mux2_1 _25163_ (.A0(_08125_),
    .A1(net2914),
    .S(_08109_),
    .X(_08126_));
 sky130_fd_sc_hd__clkbuf_1 _25164_ (.A(_08126_),
    .X(_02411_));
 sky130_fd_sc_hd__o211a_1 _25165_ (.A1(_12194_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08086_),
    .X(_08127_));
 sky130_fd_sc_hd__mux2_1 _25166_ (.A0(_08127_),
    .A1(net2563),
    .S(_08109_),
    .X(_08128_));
 sky130_fd_sc_hd__clkbuf_1 _25167_ (.A(_08128_),
    .X(_02412_));
 sky130_fd_sc_hd__o211a_1 _25168_ (.A1(_12202_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08089_),
    .X(_08129_));
 sky130_fd_sc_hd__mux2_1 _25169_ (.A0(_08129_),
    .A1(net2556),
    .S(_08109_),
    .X(_08130_));
 sky130_fd_sc_hd__clkbuf_1 _25170_ (.A(_08130_),
    .X(_02413_));
 sky130_fd_sc_hd__o211a_1 _25171_ (.A1(_12210_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08092_),
    .X(_08131_));
 sky130_fd_sc_hd__mux2_1 _25172_ (.A0(_08131_),
    .A1(net2970),
    .S(_08109_),
    .X(_08132_));
 sky130_fd_sc_hd__clkbuf_1 _25173_ (.A(_08132_),
    .X(_02414_));
 sky130_fd_sc_hd__o211a_1 _25174_ (.A1(_12218_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08095_),
    .X(_08133_));
 sky130_fd_sc_hd__mux2_1 _25175_ (.A0(_08133_),
    .A1(net2183),
    .S(_08109_),
    .X(_08134_));
 sky130_fd_sc_hd__clkbuf_1 _25176_ (.A(_08134_),
    .X(_02415_));
 sky130_fd_sc_hd__o211a_1 _25177_ (.A1(_12226_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08098_),
    .X(_08135_));
 sky130_fd_sc_hd__mux2_1 _25178_ (.A0(_08135_),
    .A1(net3191),
    .S(_08109_),
    .X(_08136_));
 sky130_fd_sc_hd__clkbuf_1 _25179_ (.A(_08136_),
    .X(_02416_));
 sky130_fd_sc_hd__o211a_1 _25180_ (.A1(_12234_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08101_),
    .X(_08137_));
 sky130_fd_sc_hd__mux2_1 _25181_ (.A0(_08137_),
    .A1(net2976),
    .S(_08109_),
    .X(_08138_));
 sky130_fd_sc_hd__clkbuf_1 _25182_ (.A(_08138_),
    .X(_02417_));
 sky130_fd_sc_hd__o211a_1 _25183_ (.A1(_12242_),
    .A2(_08082_),
    .B1(_08107_),
    .C1(_08104_),
    .X(_08139_));
 sky130_fd_sc_hd__mux2_1 _25184_ (.A0(_08139_),
    .A1(net3096),
    .S(_08109_),
    .X(_08140_));
 sky130_fd_sc_hd__clkbuf_1 _25185_ (.A(_08140_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_2 _25186_ (.A(_03371_),
    .B(_12177_),
    .Y(_08141_));
 sky130_fd_sc_hd__a21bo_1 _25187_ (.A1(_08141_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_08142_));
 sky130_fd_sc_hd__clkbuf_8 _25188_ (.A(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__mux2_1 _25189_ (.A0(_07699_),
    .A1(net2429),
    .S(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__clkbuf_1 _25190_ (.A(_08144_),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _25191_ (.A0(_07703_),
    .A1(net2851),
    .S(_08143_),
    .X(_08145_));
 sky130_fd_sc_hd__clkbuf_1 _25192_ (.A(_08145_),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _25193_ (.A0(_07705_),
    .A1(net2310),
    .S(_08143_),
    .X(_08146_));
 sky130_fd_sc_hd__clkbuf_1 _25194_ (.A(_08146_),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _25195_ (.A0(_07707_),
    .A1(net3185),
    .S(_08143_),
    .X(_08147_));
 sky130_fd_sc_hd__clkbuf_1 _25196_ (.A(_08147_),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _25197_ (.A0(_07709_),
    .A1(net2542),
    .S(_08143_),
    .X(_08148_));
 sky130_fd_sc_hd__clkbuf_1 _25198_ (.A(_08148_),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _25199_ (.A0(_07711_),
    .A1(net3690),
    .S(_08143_),
    .X(_08149_));
 sky130_fd_sc_hd__clkbuf_1 _25200_ (.A(_08149_),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _25201_ (.A0(_07713_),
    .A1(net3205),
    .S(_08143_),
    .X(_08150_));
 sky130_fd_sc_hd__clkbuf_1 _25202_ (.A(_08150_),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _25203_ (.A0(_07715_),
    .A1(net2421),
    .S(_08143_),
    .X(_08151_));
 sky130_fd_sc_hd__clkbuf_1 _25204_ (.A(_08151_),
    .X(_02426_));
 sky130_fd_sc_hd__buf_4 _25205_ (.A(_08141_),
    .X(_08152_));
 sky130_fd_sc_hd__buf_4 _25206_ (.A(_06885_),
    .X(_08153_));
 sky130_fd_sc_hd__buf_4 _25207_ (.A(_08141_),
    .X(_08154_));
 sky130_fd_sc_hd__nand2_1 _25208_ (.A(_08154_),
    .B(_12184_),
    .Y(_08155_));
 sky130_fd_sc_hd__o211a_1 _25209_ (.A1(_02850_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__mux2_1 _25210_ (.A0(_08156_),
    .A1(net3083),
    .S(_08143_),
    .X(_08157_));
 sky130_fd_sc_hd__clkbuf_1 _25211_ (.A(_08157_),
    .X(_02427_));
 sky130_fd_sc_hd__nand2_1 _25212_ (.A(_08154_),
    .B(_12197_),
    .Y(_08158_));
 sky130_fd_sc_hd__o211a_1 _25213_ (.A1(_02860_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08158_),
    .X(_08159_));
 sky130_fd_sc_hd__mux2_1 _25214_ (.A0(_08159_),
    .A1(net3731),
    .S(_08143_),
    .X(_08160_));
 sky130_fd_sc_hd__clkbuf_1 _25215_ (.A(_08160_),
    .X(_02428_));
 sky130_fd_sc_hd__nand2_1 _25216_ (.A(_08154_),
    .B(_12205_),
    .Y(_08161_));
 sky130_fd_sc_hd__o211a_1 _25217_ (.A1(_02867_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__mux2_1 _25218_ (.A0(_08162_),
    .A1(net2394),
    .S(_08143_),
    .X(_08163_));
 sky130_fd_sc_hd__clkbuf_1 _25219_ (.A(_08163_),
    .X(_02429_));
 sky130_fd_sc_hd__nand2_1 _25220_ (.A(_08154_),
    .B(_12213_),
    .Y(_08164_));
 sky130_fd_sc_hd__o211a_1 _25221_ (.A1(_02874_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__mux2_1 _25222_ (.A0(_08165_),
    .A1(net3570),
    .S(_08143_),
    .X(_08166_));
 sky130_fd_sc_hd__clkbuf_1 _25223_ (.A(_08166_),
    .X(_02430_));
 sky130_fd_sc_hd__nand2_1 _25224_ (.A(_08154_),
    .B(_12221_),
    .Y(_08167_));
 sky130_fd_sc_hd__o211a_1 _25225_ (.A1(_02881_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__mux2_1 _25226_ (.A0(_08168_),
    .A1(net2439),
    .S(_08143_),
    .X(_08169_));
 sky130_fd_sc_hd__clkbuf_1 _25227_ (.A(_08169_),
    .X(_02431_));
 sky130_fd_sc_hd__nand2_1 _25228_ (.A(_08154_),
    .B(_12229_),
    .Y(_08170_));
 sky130_fd_sc_hd__o211a_1 _25229_ (.A1(_02888_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__mux2_1 _25230_ (.A0(_08171_),
    .A1(net3740),
    .S(_08143_),
    .X(_08172_));
 sky130_fd_sc_hd__clkbuf_1 _25231_ (.A(_08172_),
    .X(_02432_));
 sky130_fd_sc_hd__nand2_1 _25232_ (.A(_08154_),
    .B(_12237_),
    .Y(_08173_));
 sky130_fd_sc_hd__o211a_1 _25233_ (.A1(_02895_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08173_),
    .X(_08174_));
 sky130_fd_sc_hd__mux2_1 _25234_ (.A0(_08174_),
    .A1(net3662),
    .S(_08143_),
    .X(_08175_));
 sky130_fd_sc_hd__clkbuf_1 _25235_ (.A(_08175_),
    .X(_02433_));
 sky130_fd_sc_hd__nand2_1 _25236_ (.A(_08154_),
    .B(_12245_),
    .Y(_08176_));
 sky130_fd_sc_hd__o211a_1 _25237_ (.A1(_02902_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__mux2_1 _25238_ (.A0(_08177_),
    .A1(net2711),
    .S(_08143_),
    .X(_08178_));
 sky130_fd_sc_hd__clkbuf_1 _25239_ (.A(_08178_),
    .X(_02434_));
 sky130_fd_sc_hd__o211a_1 _25240_ (.A1(_02910_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08155_),
    .X(_08179_));
 sky130_fd_sc_hd__clkbuf_8 _25241_ (.A(_08142_),
    .X(_08180_));
 sky130_fd_sc_hd__mux2_1 _25242_ (.A0(_08179_),
    .A1(net3477),
    .S(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__clkbuf_1 _25243_ (.A(_08181_),
    .X(_02435_));
 sky130_fd_sc_hd__o211a_1 _25244_ (.A1(_02915_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08158_),
    .X(_08182_));
 sky130_fd_sc_hd__mux2_1 _25245_ (.A0(_08182_),
    .A1(net2978),
    .S(_08180_),
    .X(_08183_));
 sky130_fd_sc_hd__clkbuf_1 _25246_ (.A(_08183_),
    .X(_02436_));
 sky130_fd_sc_hd__o211a_1 _25247_ (.A1(_02920_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08161_),
    .X(_08184_));
 sky130_fd_sc_hd__mux2_1 _25248_ (.A0(_08184_),
    .A1(net3310),
    .S(_08180_),
    .X(_08185_));
 sky130_fd_sc_hd__clkbuf_1 _25249_ (.A(_08185_),
    .X(_02437_));
 sky130_fd_sc_hd__o211a_1 _25250_ (.A1(_02926_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08164_),
    .X(_08186_));
 sky130_fd_sc_hd__mux2_1 _25251_ (.A0(_08186_),
    .A1(net2278),
    .S(_08180_),
    .X(_08187_));
 sky130_fd_sc_hd__clkbuf_1 _25252_ (.A(_08187_),
    .X(_02438_));
 sky130_fd_sc_hd__o211a_1 _25253_ (.A1(_02931_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08167_),
    .X(_08188_));
 sky130_fd_sc_hd__mux2_1 _25254_ (.A0(_08188_),
    .A1(net3340),
    .S(_08180_),
    .X(_08189_));
 sky130_fd_sc_hd__clkbuf_1 _25255_ (.A(_08189_),
    .X(_02439_));
 sky130_fd_sc_hd__o211a_1 _25256_ (.A1(_02936_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08170_),
    .X(_08190_));
 sky130_fd_sc_hd__mux2_1 _25257_ (.A0(_08190_),
    .A1(net3182),
    .S(_08180_),
    .X(_08191_));
 sky130_fd_sc_hd__clkbuf_1 _25258_ (.A(_08191_),
    .X(_02440_));
 sky130_fd_sc_hd__o211a_1 _25259_ (.A1(_02941_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08173_),
    .X(_08192_));
 sky130_fd_sc_hd__mux2_1 _25260_ (.A0(_08192_),
    .A1(net3079),
    .S(_08180_),
    .X(_08193_));
 sky130_fd_sc_hd__clkbuf_1 _25261_ (.A(_08193_),
    .X(_02441_));
 sky130_fd_sc_hd__o211a_1 _25262_ (.A1(_02946_),
    .A2(_08152_),
    .B1(_08153_),
    .C1(_08176_),
    .X(_08194_));
 sky130_fd_sc_hd__mux2_1 _25263_ (.A0(_08194_),
    .A1(net3190),
    .S(_08180_),
    .X(_08195_));
 sky130_fd_sc_hd__clkbuf_1 _25264_ (.A(_08195_),
    .X(_02442_));
 sky130_fd_sc_hd__buf_4 _25265_ (.A(_06885_),
    .X(_08196_));
 sky130_fd_sc_hd__o211a_1 _25266_ (.A1(_12169_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08155_),
    .X(_08197_));
 sky130_fd_sc_hd__mux2_1 _25267_ (.A0(_08197_),
    .A1(net2258),
    .S(_08180_),
    .X(_08198_));
 sky130_fd_sc_hd__clkbuf_1 _25268_ (.A(_08198_),
    .X(_02443_));
 sky130_fd_sc_hd__o211a_1 _25269_ (.A1(_12194_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08158_),
    .X(_08199_));
 sky130_fd_sc_hd__mux2_1 _25270_ (.A0(_08199_),
    .A1(net3261),
    .S(_08180_),
    .X(_08200_));
 sky130_fd_sc_hd__clkbuf_1 _25271_ (.A(_08200_),
    .X(_02444_));
 sky130_fd_sc_hd__o211a_1 _25272_ (.A1(_12202_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08161_),
    .X(_08201_));
 sky130_fd_sc_hd__mux2_1 _25273_ (.A0(_08201_),
    .A1(net3410),
    .S(_08180_),
    .X(_08202_));
 sky130_fd_sc_hd__clkbuf_1 _25274_ (.A(_08202_),
    .X(_02445_));
 sky130_fd_sc_hd__o211a_1 _25275_ (.A1(_12210_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08164_),
    .X(_08203_));
 sky130_fd_sc_hd__mux2_1 _25276_ (.A0(_08203_),
    .A1(net2877),
    .S(_08180_),
    .X(_08204_));
 sky130_fd_sc_hd__clkbuf_1 _25277_ (.A(_08204_),
    .X(_02446_));
 sky130_fd_sc_hd__o211a_1 _25278_ (.A1(_12218_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08167_),
    .X(_08205_));
 sky130_fd_sc_hd__mux2_1 _25279_ (.A0(_08205_),
    .A1(net3107),
    .S(_08180_),
    .X(_08206_));
 sky130_fd_sc_hd__clkbuf_1 _25280_ (.A(_08206_),
    .X(_02447_));
 sky130_fd_sc_hd__o211a_1 _25281_ (.A1(_12226_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08170_),
    .X(_08207_));
 sky130_fd_sc_hd__mux2_1 _25282_ (.A0(_08207_),
    .A1(net2655),
    .S(_08180_),
    .X(_08208_));
 sky130_fd_sc_hd__clkbuf_1 _25283_ (.A(_08208_),
    .X(_02448_));
 sky130_fd_sc_hd__o211a_1 _25284_ (.A1(_12234_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08173_),
    .X(_08209_));
 sky130_fd_sc_hd__mux2_1 _25285_ (.A0(_08209_),
    .A1(net3449),
    .S(_08180_),
    .X(_08210_));
 sky130_fd_sc_hd__clkbuf_1 _25286_ (.A(_08210_),
    .X(_02449_));
 sky130_fd_sc_hd__o211a_1 _25287_ (.A1(_12242_),
    .A2(_08154_),
    .B1(_08196_),
    .C1(_08176_),
    .X(_08211_));
 sky130_fd_sc_hd__mux2_1 _25288_ (.A0(_08211_),
    .A1(net2480),
    .S(_08180_),
    .X(_08212_));
 sky130_fd_sc_hd__clkbuf_1 _25289_ (.A(_08212_),
    .X(_02450_));
 sky130_fd_sc_hd__nand2_1 _25290_ (.A(_03443_),
    .B(_12177_),
    .Y(_08213_));
 sky130_fd_sc_hd__a21bo_1 _25291_ (.A1(_08213_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_08214_));
 sky130_fd_sc_hd__clkbuf_8 _25292_ (.A(_08214_),
    .X(_08215_));
 sky130_fd_sc_hd__mux2_1 _25293_ (.A0(_07699_),
    .A1(net2493),
    .S(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__clkbuf_1 _25294_ (.A(_08216_),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _25295_ (.A0(_07703_),
    .A1(net2945),
    .S(_08215_),
    .X(_08217_));
 sky130_fd_sc_hd__clkbuf_1 _25296_ (.A(_08217_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _25297_ (.A0(_07705_),
    .A1(net2203),
    .S(_08215_),
    .X(_08218_));
 sky130_fd_sc_hd__clkbuf_1 _25298_ (.A(_08218_),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _25299_ (.A0(_07707_),
    .A1(net2297),
    .S(_08215_),
    .X(_08219_));
 sky130_fd_sc_hd__clkbuf_1 _25300_ (.A(_08219_),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _25301_ (.A0(_07709_),
    .A1(net2231),
    .S(_08215_),
    .X(_08220_));
 sky130_fd_sc_hd__clkbuf_1 _25302_ (.A(_08220_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _25303_ (.A0(_07711_),
    .A1(net2245),
    .S(_08215_),
    .X(_08221_));
 sky130_fd_sc_hd__clkbuf_1 _25304_ (.A(_08221_),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _25305_ (.A0(_07713_),
    .A1(net3313),
    .S(_08215_),
    .X(_08222_));
 sky130_fd_sc_hd__clkbuf_1 _25306_ (.A(_08222_),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _25307_ (.A0(_07715_),
    .A1(net3131),
    .S(_08215_),
    .X(_08223_));
 sky130_fd_sc_hd__clkbuf_1 _25308_ (.A(_08223_),
    .X(_02458_));
 sky130_fd_sc_hd__buf_4 _25309_ (.A(_08213_),
    .X(_08224_));
 sky130_fd_sc_hd__buf_4 _25310_ (.A(_08213_),
    .X(_08225_));
 sky130_fd_sc_hd__nand2_1 _25311_ (.A(_08225_),
    .B(_12184_),
    .Y(_08226_));
 sky130_fd_sc_hd__o211a_1 _25312_ (.A1(_02850_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__mux2_1 _25313_ (.A0(_08227_),
    .A1(net2967),
    .S(_08215_),
    .X(_08228_));
 sky130_fd_sc_hd__clkbuf_1 _25314_ (.A(_08228_),
    .X(_02459_));
 sky130_fd_sc_hd__nand2_1 _25315_ (.A(_08225_),
    .B(_12197_),
    .Y(_08229_));
 sky130_fd_sc_hd__o211a_1 _25316_ (.A1(_02860_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__mux2_1 _25317_ (.A0(_08230_),
    .A1(net3632),
    .S(_08215_),
    .X(_08231_));
 sky130_fd_sc_hd__clkbuf_1 _25318_ (.A(_08231_),
    .X(_02460_));
 sky130_fd_sc_hd__nand2_1 _25319_ (.A(_08225_),
    .B(_12205_),
    .Y(_08232_));
 sky130_fd_sc_hd__o211a_1 _25320_ (.A1(_02867_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__mux2_1 _25321_ (.A0(_08233_),
    .A1(net3295),
    .S(_08215_),
    .X(_08234_));
 sky130_fd_sc_hd__clkbuf_1 _25322_ (.A(_08234_),
    .X(_02461_));
 sky130_fd_sc_hd__nand2_1 _25323_ (.A(_08225_),
    .B(_12213_),
    .Y(_08235_));
 sky130_fd_sc_hd__o211a_1 _25324_ (.A1(_02874_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__mux2_1 _25325_ (.A0(_08236_),
    .A1(net3063),
    .S(_08215_),
    .X(_08237_));
 sky130_fd_sc_hd__clkbuf_1 _25326_ (.A(_08237_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2_1 _25327_ (.A(_08225_),
    .B(_12221_),
    .Y(_08238_));
 sky130_fd_sc_hd__o211a_1 _25328_ (.A1(_02881_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__mux2_1 _25329_ (.A0(_08239_),
    .A1(net2608),
    .S(_08215_),
    .X(_08240_));
 sky130_fd_sc_hd__clkbuf_1 _25330_ (.A(_08240_),
    .X(_02463_));
 sky130_fd_sc_hd__nand2_1 _25331_ (.A(_08225_),
    .B(_12229_),
    .Y(_08241_));
 sky130_fd_sc_hd__o211a_1 _25332_ (.A1(_02888_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__mux2_1 _25333_ (.A0(_08242_),
    .A1(net2580),
    .S(_08215_),
    .X(_08243_));
 sky130_fd_sc_hd__clkbuf_1 _25334_ (.A(_08243_),
    .X(_02464_));
 sky130_fd_sc_hd__nand2_1 _25335_ (.A(_08225_),
    .B(_12237_),
    .Y(_08244_));
 sky130_fd_sc_hd__o211a_1 _25336_ (.A1(_02895_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__mux2_1 _25337_ (.A0(_08245_),
    .A1(net3455),
    .S(_08215_),
    .X(_08246_));
 sky130_fd_sc_hd__clkbuf_1 _25338_ (.A(_08246_),
    .X(_02465_));
 sky130_fd_sc_hd__nand2_1 _25339_ (.A(_08225_),
    .B(_12245_),
    .Y(_08247_));
 sky130_fd_sc_hd__o211a_1 _25340_ (.A1(_02902_),
    .A2(_08224_),
    .B1(_08196_),
    .C1(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__mux2_1 _25341_ (.A0(_08248_),
    .A1(net3691),
    .S(_08215_),
    .X(_08249_));
 sky130_fd_sc_hd__clkbuf_1 _25342_ (.A(_08249_),
    .X(_02466_));
 sky130_fd_sc_hd__buf_4 _25343_ (.A(_06885_),
    .X(_08250_));
 sky130_fd_sc_hd__o211a_1 _25344_ (.A1(_02910_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08226_),
    .X(_08251_));
 sky130_fd_sc_hd__clkbuf_8 _25345_ (.A(_08214_),
    .X(_08252_));
 sky130_fd_sc_hd__mux2_1 _25346_ (.A0(_08251_),
    .A1(net3831),
    .S(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__clkbuf_1 _25347_ (.A(_08253_),
    .X(_02467_));
 sky130_fd_sc_hd__o211a_1 _25348_ (.A1(_02915_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08229_),
    .X(_08254_));
 sky130_fd_sc_hd__mux2_1 _25349_ (.A0(_08254_),
    .A1(net3338),
    .S(_08252_),
    .X(_08255_));
 sky130_fd_sc_hd__clkbuf_1 _25350_ (.A(_08255_),
    .X(_02468_));
 sky130_fd_sc_hd__o211a_1 _25351_ (.A1(_02920_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08232_),
    .X(_08256_));
 sky130_fd_sc_hd__mux2_1 _25352_ (.A0(_08256_),
    .A1(net3858),
    .S(_08252_),
    .X(_08257_));
 sky130_fd_sc_hd__clkbuf_1 _25353_ (.A(_08257_),
    .X(_02469_));
 sky130_fd_sc_hd__o211a_1 _25354_ (.A1(_02926_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08235_),
    .X(_08258_));
 sky130_fd_sc_hd__mux2_1 _25355_ (.A0(_08258_),
    .A1(net3664),
    .S(_08252_),
    .X(_08259_));
 sky130_fd_sc_hd__clkbuf_1 _25356_ (.A(_08259_),
    .X(_02470_));
 sky130_fd_sc_hd__o211a_1 _25357_ (.A1(_02931_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08238_),
    .X(_08260_));
 sky130_fd_sc_hd__mux2_1 _25358_ (.A0(_08260_),
    .A1(net3349),
    .S(_08252_),
    .X(_08261_));
 sky130_fd_sc_hd__clkbuf_1 _25359_ (.A(_08261_),
    .X(_02471_));
 sky130_fd_sc_hd__o211a_1 _25360_ (.A1(_02936_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08241_),
    .X(_08262_));
 sky130_fd_sc_hd__mux2_1 _25361_ (.A0(_08262_),
    .A1(net3709),
    .S(_08252_),
    .X(_08263_));
 sky130_fd_sc_hd__clkbuf_1 _25362_ (.A(_08263_),
    .X(_02472_));
 sky130_fd_sc_hd__o211a_1 _25363_ (.A1(_02941_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08244_),
    .X(_08264_));
 sky130_fd_sc_hd__mux2_1 _25364_ (.A0(_08264_),
    .A1(net3775),
    .S(_08252_),
    .X(_08265_));
 sky130_fd_sc_hd__clkbuf_1 _25365_ (.A(_08265_),
    .X(_02473_));
 sky130_fd_sc_hd__o211a_1 _25366_ (.A1(_02946_),
    .A2(_08224_),
    .B1(_08250_),
    .C1(_08247_),
    .X(_08266_));
 sky130_fd_sc_hd__mux2_1 _25367_ (.A0(_08266_),
    .A1(net3859),
    .S(_08252_),
    .X(_08267_));
 sky130_fd_sc_hd__clkbuf_1 _25368_ (.A(_08267_),
    .X(_02474_));
 sky130_fd_sc_hd__o211a_1 _25369_ (.A1(_12169_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08226_),
    .X(_08268_));
 sky130_fd_sc_hd__mux2_1 _25370_ (.A0(_08268_),
    .A1(net3930),
    .S(_08252_),
    .X(_08269_));
 sky130_fd_sc_hd__clkbuf_1 _25371_ (.A(_08269_),
    .X(_02475_));
 sky130_fd_sc_hd__o211a_1 _25372_ (.A1(_12194_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08229_),
    .X(_08270_));
 sky130_fd_sc_hd__mux2_1 _25373_ (.A0(_08270_),
    .A1(net3925),
    .S(_08252_),
    .X(_08271_));
 sky130_fd_sc_hd__clkbuf_1 _25374_ (.A(_08271_),
    .X(_02476_));
 sky130_fd_sc_hd__o211a_1 _25375_ (.A1(_12202_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08232_),
    .X(_08272_));
 sky130_fd_sc_hd__mux2_1 _25376_ (.A0(_08272_),
    .A1(net3924),
    .S(_08252_),
    .X(_08273_));
 sky130_fd_sc_hd__clkbuf_1 _25377_ (.A(_08273_),
    .X(_02477_));
 sky130_fd_sc_hd__o211a_1 _25378_ (.A1(_12210_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08235_),
    .X(_08274_));
 sky130_fd_sc_hd__mux2_1 _25379_ (.A0(_08274_),
    .A1(net3883),
    .S(_08252_),
    .X(_08275_));
 sky130_fd_sc_hd__clkbuf_1 _25380_ (.A(_08275_),
    .X(_02478_));
 sky130_fd_sc_hd__o211a_1 _25381_ (.A1(_12218_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08238_),
    .X(_08276_));
 sky130_fd_sc_hd__mux2_1 _25382_ (.A0(_08276_),
    .A1(net3919),
    .S(_08252_),
    .X(_08277_));
 sky130_fd_sc_hd__clkbuf_1 _25383_ (.A(_08277_),
    .X(_02479_));
 sky130_fd_sc_hd__o211a_1 _25384_ (.A1(_12226_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08241_),
    .X(_08278_));
 sky130_fd_sc_hd__mux2_1 _25385_ (.A0(_08278_),
    .A1(net3909),
    .S(_08252_),
    .X(_08279_));
 sky130_fd_sc_hd__clkbuf_1 _25386_ (.A(_08279_),
    .X(_02480_));
 sky130_fd_sc_hd__o211a_1 _25387_ (.A1(_12234_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08244_),
    .X(_08280_));
 sky130_fd_sc_hd__mux2_1 _25388_ (.A0(_08280_),
    .A1(net3920),
    .S(_08252_),
    .X(_08281_));
 sky130_fd_sc_hd__clkbuf_1 _25389_ (.A(_08281_),
    .X(_02481_));
 sky130_fd_sc_hd__o211a_1 _25390_ (.A1(_12242_),
    .A2(_08225_),
    .B1(_08250_),
    .C1(_08247_),
    .X(_08282_));
 sky130_fd_sc_hd__mux2_1 _25391_ (.A0(_08282_),
    .A1(net3917),
    .S(_08252_),
    .X(_08283_));
 sky130_fd_sc_hd__clkbuf_1 _25392_ (.A(_08283_),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_2 _25393_ (.A(_03519_),
    .B(_12177_),
    .Y(_08284_));
 sky130_fd_sc_hd__a21bo_1 _25394_ (.A1(_08284_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_08285_));
 sky130_fd_sc_hd__buf_6 _25395_ (.A(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__mux2_1 _25396_ (.A0(_07699_),
    .A1(net2286),
    .S(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__clkbuf_1 _25397_ (.A(_08287_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _25398_ (.A0(_07703_),
    .A1(net2621),
    .S(_08286_),
    .X(_08288_));
 sky130_fd_sc_hd__clkbuf_1 _25399_ (.A(_08288_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _25400_ (.A0(_07705_),
    .A1(net2471),
    .S(_08286_),
    .X(_08289_));
 sky130_fd_sc_hd__clkbuf_1 _25401_ (.A(_08289_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _25402_ (.A0(_07707_),
    .A1(net3080),
    .S(_08286_),
    .X(_08290_));
 sky130_fd_sc_hd__clkbuf_1 _25403_ (.A(_08290_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _25404_ (.A0(_07709_),
    .A1(net2350),
    .S(_08286_),
    .X(_08291_));
 sky130_fd_sc_hd__clkbuf_1 _25405_ (.A(_08291_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _25406_ (.A0(_07711_),
    .A1(net2968),
    .S(_08286_),
    .X(_08292_));
 sky130_fd_sc_hd__clkbuf_1 _25407_ (.A(_08292_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _25408_ (.A0(_07713_),
    .A1(net2279),
    .S(_08286_),
    .X(_08293_));
 sky130_fd_sc_hd__clkbuf_1 _25409_ (.A(_08293_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _25410_ (.A0(_07715_),
    .A1(net3249),
    .S(_08286_),
    .X(_08294_));
 sky130_fd_sc_hd__clkbuf_1 _25411_ (.A(_08294_),
    .X(_02490_));
 sky130_fd_sc_hd__buf_4 _25412_ (.A(_08284_),
    .X(_08295_));
 sky130_fd_sc_hd__buf_4 _25413_ (.A(_06885_),
    .X(_08296_));
 sky130_fd_sc_hd__buf_4 _25414_ (.A(_08284_),
    .X(_08297_));
 sky130_fd_sc_hd__nand2_1 _25415_ (.A(_08297_),
    .B(_12184_),
    .Y(_08298_));
 sky130_fd_sc_hd__o211a_1 _25416_ (.A1(_02850_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__mux2_1 _25417_ (.A0(_08299_),
    .A1(net2665),
    .S(_08286_),
    .X(_08300_));
 sky130_fd_sc_hd__clkbuf_1 _25418_ (.A(_08300_),
    .X(_02491_));
 sky130_fd_sc_hd__nand2_1 _25419_ (.A(_08297_),
    .B(_12197_),
    .Y(_08301_));
 sky130_fd_sc_hd__o211a_1 _25420_ (.A1(_02860_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__mux2_1 _25421_ (.A0(_08302_),
    .A1(net2979),
    .S(_08286_),
    .X(_08303_));
 sky130_fd_sc_hd__clkbuf_1 _25422_ (.A(_08303_),
    .X(_02492_));
 sky130_fd_sc_hd__nand2_1 _25423_ (.A(_08297_),
    .B(_12205_),
    .Y(_08304_));
 sky130_fd_sc_hd__o211a_1 _25424_ (.A1(_02867_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__mux2_1 _25425_ (.A0(_08305_),
    .A1(net2805),
    .S(_08286_),
    .X(_08306_));
 sky130_fd_sc_hd__clkbuf_1 _25426_ (.A(_08306_),
    .X(_02493_));
 sky130_fd_sc_hd__nand2_1 _25427_ (.A(_08297_),
    .B(_12213_),
    .Y(_08307_));
 sky130_fd_sc_hd__o211a_1 _25428_ (.A1(_02874_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__mux2_1 _25429_ (.A0(_08308_),
    .A1(net2881),
    .S(_08286_),
    .X(_08309_));
 sky130_fd_sc_hd__clkbuf_1 _25430_ (.A(_08309_),
    .X(_02494_));
 sky130_fd_sc_hd__nand2_1 _25431_ (.A(_08297_),
    .B(_12221_),
    .Y(_08310_));
 sky130_fd_sc_hd__o211a_1 _25432_ (.A1(_02881_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08310_),
    .X(_08311_));
 sky130_fd_sc_hd__mux2_1 _25433_ (.A0(_08311_),
    .A1(net2952),
    .S(_08286_),
    .X(_08312_));
 sky130_fd_sc_hd__clkbuf_1 _25434_ (.A(_08312_),
    .X(_02495_));
 sky130_fd_sc_hd__nand2_1 _25435_ (.A(_08297_),
    .B(_12229_),
    .Y(_08313_));
 sky130_fd_sc_hd__o211a_1 _25436_ (.A1(_02888_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__mux2_1 _25437_ (.A0(_08314_),
    .A1(net2640),
    .S(_08286_),
    .X(_08315_));
 sky130_fd_sc_hd__clkbuf_1 _25438_ (.A(_08315_),
    .X(_02496_));
 sky130_fd_sc_hd__nand2_1 _25439_ (.A(_08297_),
    .B(_12237_),
    .Y(_08316_));
 sky130_fd_sc_hd__o211a_1 _25440_ (.A1(_02895_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__mux2_1 _25441_ (.A0(_08317_),
    .A1(net2925),
    .S(_08286_),
    .X(_08318_));
 sky130_fd_sc_hd__clkbuf_1 _25442_ (.A(_08318_),
    .X(_02497_));
 sky130_fd_sc_hd__nand2_1 _25443_ (.A(_08297_),
    .B(_12245_),
    .Y(_08319_));
 sky130_fd_sc_hd__o211a_1 _25444_ (.A1(_02902_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__mux2_1 _25445_ (.A0(_08320_),
    .A1(net2998),
    .S(_08286_),
    .X(_08321_));
 sky130_fd_sc_hd__clkbuf_1 _25446_ (.A(_08321_),
    .X(_02498_));
 sky130_fd_sc_hd__o211a_1 _25447_ (.A1(_02910_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08298_),
    .X(_08322_));
 sky130_fd_sc_hd__clkbuf_8 _25448_ (.A(_08285_),
    .X(_08323_));
 sky130_fd_sc_hd__mux2_1 _25449_ (.A0(_08322_),
    .A1(net3454),
    .S(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__clkbuf_1 _25450_ (.A(_08324_),
    .X(_02499_));
 sky130_fd_sc_hd__o211a_1 _25451_ (.A1(_02915_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08301_),
    .X(_08325_));
 sky130_fd_sc_hd__mux2_1 _25452_ (.A0(_08325_),
    .A1(net2762),
    .S(_08323_),
    .X(_08326_));
 sky130_fd_sc_hd__clkbuf_1 _25453_ (.A(_08326_),
    .X(_02500_));
 sky130_fd_sc_hd__o211a_1 _25454_ (.A1(_02920_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08304_),
    .X(_08327_));
 sky130_fd_sc_hd__mux2_1 _25455_ (.A0(_08327_),
    .A1(net2333),
    .S(_08323_),
    .X(_08328_));
 sky130_fd_sc_hd__clkbuf_1 _25456_ (.A(_08328_),
    .X(_02501_));
 sky130_fd_sc_hd__o211a_1 _25457_ (.A1(_02926_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08307_),
    .X(_08329_));
 sky130_fd_sc_hd__mux2_1 _25458_ (.A0(_08329_),
    .A1(net3534),
    .S(_08323_),
    .X(_08330_));
 sky130_fd_sc_hd__clkbuf_1 _25459_ (.A(_08330_),
    .X(_02502_));
 sky130_fd_sc_hd__o211a_1 _25460_ (.A1(_02931_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08310_),
    .X(_08331_));
 sky130_fd_sc_hd__mux2_1 _25461_ (.A0(_08331_),
    .A1(net3105),
    .S(_08323_),
    .X(_08332_));
 sky130_fd_sc_hd__clkbuf_1 _25462_ (.A(_08332_),
    .X(_02503_));
 sky130_fd_sc_hd__o211a_1 _25463_ (.A1(_02936_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08313_),
    .X(_08333_));
 sky130_fd_sc_hd__mux2_1 _25464_ (.A0(_08333_),
    .A1(net3002),
    .S(_08323_),
    .X(_08334_));
 sky130_fd_sc_hd__clkbuf_1 _25465_ (.A(_08334_),
    .X(_02504_));
 sky130_fd_sc_hd__o211a_1 _25466_ (.A1(_02941_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08316_),
    .X(_08335_));
 sky130_fd_sc_hd__mux2_1 _25467_ (.A0(_08335_),
    .A1(net3431),
    .S(_08323_),
    .X(_08336_));
 sky130_fd_sc_hd__clkbuf_1 _25468_ (.A(_08336_),
    .X(_02505_));
 sky130_fd_sc_hd__o211a_1 _25469_ (.A1(_02946_),
    .A2(_08295_),
    .B1(_08296_),
    .C1(_08319_),
    .X(_08337_));
 sky130_fd_sc_hd__mux2_1 _25470_ (.A0(_08337_),
    .A1(net2632),
    .S(_08323_),
    .X(_08338_));
 sky130_fd_sc_hd__clkbuf_1 _25471_ (.A(_08338_),
    .X(_02506_));
 sky130_fd_sc_hd__buf_4 _25472_ (.A(_06885_),
    .X(_08339_));
 sky130_fd_sc_hd__o211a_1 _25473_ (.A1(_12169_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08298_),
    .X(_08340_));
 sky130_fd_sc_hd__mux2_1 _25474_ (.A0(_08340_),
    .A1(net2657),
    .S(_08323_),
    .X(_08341_));
 sky130_fd_sc_hd__clkbuf_1 _25475_ (.A(_08341_),
    .X(_02507_));
 sky130_fd_sc_hd__o211a_1 _25476_ (.A1(_12194_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08301_),
    .X(_08342_));
 sky130_fd_sc_hd__mux2_1 _25477_ (.A0(_08342_),
    .A1(net3161),
    .S(_08323_),
    .X(_08343_));
 sky130_fd_sc_hd__clkbuf_1 _25478_ (.A(_08343_),
    .X(_02508_));
 sky130_fd_sc_hd__o211a_1 _25479_ (.A1(_12202_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08304_),
    .X(_08344_));
 sky130_fd_sc_hd__mux2_1 _25480_ (.A0(_08344_),
    .A1(net2950),
    .S(_08323_),
    .X(_08345_));
 sky130_fd_sc_hd__clkbuf_1 _25481_ (.A(_08345_),
    .X(_02509_));
 sky130_fd_sc_hd__o211a_1 _25482_ (.A1(_12210_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08307_),
    .X(_08346_));
 sky130_fd_sc_hd__mux2_1 _25483_ (.A0(_08346_),
    .A1(net3332),
    .S(_08323_),
    .X(_08347_));
 sky130_fd_sc_hd__clkbuf_1 _25484_ (.A(_08347_),
    .X(_02510_));
 sky130_fd_sc_hd__o211a_1 _25485_ (.A1(_12218_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08310_),
    .X(_08348_));
 sky130_fd_sc_hd__mux2_1 _25486_ (.A0(_08348_),
    .A1(net2329),
    .S(_08323_),
    .X(_08349_));
 sky130_fd_sc_hd__clkbuf_1 _25487_ (.A(_08349_),
    .X(_02511_));
 sky130_fd_sc_hd__o211a_1 _25488_ (.A1(_12226_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08313_),
    .X(_08350_));
 sky130_fd_sc_hd__mux2_1 _25489_ (.A0(_08350_),
    .A1(net2889),
    .S(_08323_),
    .X(_08351_));
 sky130_fd_sc_hd__clkbuf_1 _25490_ (.A(_08351_),
    .X(_02512_));
 sky130_fd_sc_hd__o211a_1 _25491_ (.A1(_12234_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08316_),
    .X(_08352_));
 sky130_fd_sc_hd__mux2_1 _25492_ (.A0(_08352_),
    .A1(net2516),
    .S(_08323_),
    .X(_08353_));
 sky130_fd_sc_hd__clkbuf_1 _25493_ (.A(_08353_),
    .X(_02513_));
 sky130_fd_sc_hd__o211a_1 _25494_ (.A1(_12242_),
    .A2(_08297_),
    .B1(_08339_),
    .C1(_08319_),
    .X(_08354_));
 sky130_fd_sc_hd__mux2_1 _25495_ (.A0(_08354_),
    .A1(net2483),
    .S(_08323_),
    .X(_08355_));
 sky130_fd_sc_hd__clkbuf_1 _25496_ (.A(_08355_),
    .X(_02514_));
 sky130_fd_sc_hd__nand2_2 _25497_ (.A(_03591_),
    .B(_12177_),
    .Y(_08356_));
 sky130_fd_sc_hd__a21bo_1 _25498_ (.A1(_08356_),
    .A2(_06534_),
    .B1_N(_06384_),
    .X(_08357_));
 sky130_fd_sc_hd__clkbuf_8 _25499_ (.A(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__mux2_1 _25500_ (.A0(_07699_),
    .A1(net2202),
    .S(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__clkbuf_1 _25501_ (.A(_08359_),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _25502_ (.A0(_07703_),
    .A1(net2478),
    .S(_08358_),
    .X(_08360_));
 sky130_fd_sc_hd__clkbuf_1 _25503_ (.A(_08360_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _25504_ (.A0(_07705_),
    .A1(net2253),
    .S(_08358_),
    .X(_08361_));
 sky130_fd_sc_hd__clkbuf_1 _25505_ (.A(_08361_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _25506_ (.A0(_07707_),
    .A1(net3571),
    .S(_08358_),
    .X(_08362_));
 sky130_fd_sc_hd__clkbuf_1 _25507_ (.A(_08362_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _25508_ (.A0(_07709_),
    .A1(net3011),
    .S(_08358_),
    .X(_08363_));
 sky130_fd_sc_hd__clkbuf_1 _25509_ (.A(_08363_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _25510_ (.A0(_07711_),
    .A1(net2863),
    .S(_08358_),
    .X(_08364_));
 sky130_fd_sc_hd__clkbuf_1 _25511_ (.A(_08364_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _25512_ (.A0(_07713_),
    .A1(net2247),
    .S(_08358_),
    .X(_08365_));
 sky130_fd_sc_hd__clkbuf_1 _25513_ (.A(_08365_),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _25514_ (.A0(_07715_),
    .A1(net2307),
    .S(_08358_),
    .X(_08366_));
 sky130_fd_sc_hd__clkbuf_1 _25515_ (.A(_08366_),
    .X(_02522_));
 sky130_fd_sc_hd__buf_4 _25516_ (.A(_08356_),
    .X(_08367_));
 sky130_fd_sc_hd__buf_4 _25517_ (.A(_08356_),
    .X(_08368_));
 sky130_fd_sc_hd__nand2_1 _25518_ (.A(_08368_),
    .B(_12184_),
    .Y(_08369_));
 sky130_fd_sc_hd__o211a_1 _25519_ (.A1(_02850_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08369_),
    .X(_08370_));
 sky130_fd_sc_hd__mux2_1 _25520_ (.A0(_08370_),
    .A1(net3305),
    .S(_08358_),
    .X(_08371_));
 sky130_fd_sc_hd__clkbuf_1 _25521_ (.A(_08371_),
    .X(_02523_));
 sky130_fd_sc_hd__nand2_1 _25522_ (.A(_08368_),
    .B(_12197_),
    .Y(_08372_));
 sky130_fd_sc_hd__o211a_1 _25523_ (.A1(_02860_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__mux2_1 _25524_ (.A0(_08373_),
    .A1(net3257),
    .S(_08358_),
    .X(_08374_));
 sky130_fd_sc_hd__clkbuf_1 _25525_ (.A(_08374_),
    .X(_02524_));
 sky130_fd_sc_hd__nand2_1 _25526_ (.A(_08368_),
    .B(_12205_),
    .Y(_08375_));
 sky130_fd_sc_hd__o211a_1 _25527_ (.A1(_02867_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__mux2_1 _25528_ (.A0(_08376_),
    .A1(net3466),
    .S(_08358_),
    .X(_08377_));
 sky130_fd_sc_hd__clkbuf_1 _25529_ (.A(_08377_),
    .X(_02525_));
 sky130_fd_sc_hd__nand2_1 _25530_ (.A(_08368_),
    .B(_12213_),
    .Y(_08378_));
 sky130_fd_sc_hd__o211a_1 _25531_ (.A1(_02874_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__mux2_1 _25532_ (.A0(_08379_),
    .A1(net2857),
    .S(_08358_),
    .X(_08380_));
 sky130_fd_sc_hd__clkbuf_1 _25533_ (.A(_08380_),
    .X(_02526_));
 sky130_fd_sc_hd__nand2_1 _25534_ (.A(_08368_),
    .B(_12221_),
    .Y(_08381_));
 sky130_fd_sc_hd__o211a_1 _25535_ (.A1(_02881_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__mux2_1 _25536_ (.A0(_08382_),
    .A1(net2984),
    .S(_08358_),
    .X(_08383_));
 sky130_fd_sc_hd__clkbuf_1 _25537_ (.A(_08383_),
    .X(_02527_));
 sky130_fd_sc_hd__nand2_1 _25538_ (.A(_08368_),
    .B(_12229_),
    .Y(_08384_));
 sky130_fd_sc_hd__o211a_1 _25539_ (.A1(_02888_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__mux2_1 _25540_ (.A0(_08385_),
    .A1(net3353),
    .S(_08358_),
    .X(_08386_));
 sky130_fd_sc_hd__clkbuf_1 _25541_ (.A(_08386_),
    .X(_02528_));
 sky130_fd_sc_hd__nand2_1 _25542_ (.A(_08368_),
    .B(_12237_),
    .Y(_08387_));
 sky130_fd_sc_hd__o211a_1 _25543_ (.A1(_02895_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__mux2_1 _25544_ (.A0(_08388_),
    .A1(net3169),
    .S(_08358_),
    .X(_08389_));
 sky130_fd_sc_hd__clkbuf_1 _25545_ (.A(_08389_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _25546_ (.A(_08368_),
    .B(_12245_),
    .Y(_08390_));
 sky130_fd_sc_hd__o211a_1 _25547_ (.A1(_02902_),
    .A2(_08367_),
    .B1(_08339_),
    .C1(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__mux2_1 _25548_ (.A0(_08391_),
    .A1(net2567),
    .S(_08358_),
    .X(_08392_));
 sky130_fd_sc_hd__clkbuf_1 _25549_ (.A(_08392_),
    .X(_02530_));
 sky130_fd_sc_hd__buf_4 _25550_ (.A(_09125_),
    .X(_08393_));
 sky130_fd_sc_hd__o211a_1 _25551_ (.A1(_02910_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08369_),
    .X(_08394_));
 sky130_fd_sc_hd__clkbuf_8 _25552_ (.A(_08357_),
    .X(_08395_));
 sky130_fd_sc_hd__mux2_1 _25553_ (.A0(_08394_),
    .A1(net3291),
    .S(_08395_),
    .X(_08396_));
 sky130_fd_sc_hd__clkbuf_1 _25554_ (.A(_08396_),
    .X(_02531_));
 sky130_fd_sc_hd__o211a_1 _25555_ (.A1(_02915_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08372_),
    .X(_08397_));
 sky130_fd_sc_hd__mux2_1 _25556_ (.A0(_08397_),
    .A1(net3104),
    .S(_08395_),
    .X(_08398_));
 sky130_fd_sc_hd__clkbuf_1 _25557_ (.A(_08398_),
    .X(_02532_));
 sky130_fd_sc_hd__o211a_1 _25558_ (.A1(_02920_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08375_),
    .X(_08399_));
 sky130_fd_sc_hd__mux2_1 _25559_ (.A0(_08399_),
    .A1(net3342),
    .S(_08395_),
    .X(_08400_));
 sky130_fd_sc_hd__clkbuf_1 _25560_ (.A(_08400_),
    .X(_02533_));
 sky130_fd_sc_hd__o211a_1 _25561_ (.A1(_02926_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08378_),
    .X(_08401_));
 sky130_fd_sc_hd__mux2_1 _25562_ (.A0(_08401_),
    .A1(net2955),
    .S(_08395_),
    .X(_08402_));
 sky130_fd_sc_hd__clkbuf_1 _25563_ (.A(_08402_),
    .X(_02534_));
 sky130_fd_sc_hd__o211a_1 _25564_ (.A1(_02931_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08381_),
    .X(_08403_));
 sky130_fd_sc_hd__mux2_1 _25565_ (.A0(_08403_),
    .A1(net3329),
    .S(_08395_),
    .X(_08404_));
 sky130_fd_sc_hd__clkbuf_1 _25566_ (.A(_08404_),
    .X(_02535_));
 sky130_fd_sc_hd__o211a_1 _25567_ (.A1(_02936_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08384_),
    .X(_08405_));
 sky130_fd_sc_hd__mux2_1 _25568_ (.A0(_08405_),
    .A1(net2739),
    .S(_08395_),
    .X(_08406_));
 sky130_fd_sc_hd__clkbuf_1 _25569_ (.A(_08406_),
    .X(_02536_));
 sky130_fd_sc_hd__o211a_1 _25570_ (.A1(_02941_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08387_),
    .X(_08407_));
 sky130_fd_sc_hd__mux2_1 _25571_ (.A0(_08407_),
    .A1(net2742),
    .S(_08395_),
    .X(_08408_));
 sky130_fd_sc_hd__clkbuf_1 _25572_ (.A(_08408_),
    .X(_02537_));
 sky130_fd_sc_hd__o211a_1 _25573_ (.A1(_02946_),
    .A2(_08367_),
    .B1(_08393_),
    .C1(_08390_),
    .X(_08409_));
 sky130_fd_sc_hd__mux2_1 _25574_ (.A0(_08409_),
    .A1(net3087),
    .S(_08395_),
    .X(_08410_));
 sky130_fd_sc_hd__clkbuf_1 _25575_ (.A(_08410_),
    .X(_02538_));
 sky130_fd_sc_hd__o211a_1 _25576_ (.A1(_12169_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08369_),
    .X(_08411_));
 sky130_fd_sc_hd__mux2_1 _25577_ (.A0(_08411_),
    .A1(net2551),
    .S(_08395_),
    .X(_08412_));
 sky130_fd_sc_hd__clkbuf_1 _25578_ (.A(_08412_),
    .X(_02539_));
 sky130_fd_sc_hd__o211a_1 _25579_ (.A1(_12194_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08372_),
    .X(_08413_));
 sky130_fd_sc_hd__mux2_1 _25580_ (.A0(_08413_),
    .A1(net2935),
    .S(_08395_),
    .X(_08414_));
 sky130_fd_sc_hd__clkbuf_1 _25581_ (.A(_08414_),
    .X(_02540_));
 sky130_fd_sc_hd__o211a_1 _25582_ (.A1(_12202_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08375_),
    .X(_08415_));
 sky130_fd_sc_hd__mux2_1 _25583_ (.A0(_08415_),
    .A1(net2555),
    .S(_08395_),
    .X(_08416_));
 sky130_fd_sc_hd__clkbuf_1 _25584_ (.A(_08416_),
    .X(_02541_));
 sky130_fd_sc_hd__o211a_1 _25585_ (.A1(_12210_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08378_),
    .X(_08417_));
 sky130_fd_sc_hd__mux2_1 _25586_ (.A0(_08417_),
    .A1(net3546),
    .S(_08395_),
    .X(_08418_));
 sky130_fd_sc_hd__clkbuf_1 _25587_ (.A(_08418_),
    .X(_02542_));
 sky130_fd_sc_hd__o211a_1 _25588_ (.A1(_12218_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08381_),
    .X(_08419_));
 sky130_fd_sc_hd__mux2_1 _25589_ (.A0(_08419_),
    .A1(net3542),
    .S(_08395_),
    .X(_08420_));
 sky130_fd_sc_hd__clkbuf_1 _25590_ (.A(_08420_),
    .X(_02543_));
 sky130_fd_sc_hd__o211a_1 _25591_ (.A1(_12226_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08384_),
    .X(_08421_));
 sky130_fd_sc_hd__mux2_1 _25592_ (.A0(_08421_),
    .A1(net3553),
    .S(_08395_),
    .X(_08422_));
 sky130_fd_sc_hd__clkbuf_1 _25593_ (.A(_08422_),
    .X(_02544_));
 sky130_fd_sc_hd__o211a_1 _25594_ (.A1(_12234_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08387_),
    .X(_08423_));
 sky130_fd_sc_hd__mux2_1 _25595_ (.A0(_08423_),
    .A1(net2449),
    .S(_08395_),
    .X(_08424_));
 sky130_fd_sc_hd__clkbuf_1 _25596_ (.A(_08424_),
    .X(_02545_));
 sky130_fd_sc_hd__o211a_1 _25597_ (.A1(_12242_),
    .A2(_08368_),
    .B1(_08393_),
    .C1(_08390_),
    .X(_08425_));
 sky130_fd_sc_hd__mux2_1 _25598_ (.A0(_08425_),
    .A1(net2553),
    .S(_08395_),
    .X(_08426_));
 sky130_fd_sc_hd__clkbuf_1 _25599_ (.A(_08426_),
    .X(_02546_));
 sky130_fd_sc_hd__nand2_1 _25600_ (.A(_03664_),
    .B(_12177_),
    .Y(_08427_));
 sky130_fd_sc_hd__a21bo_1 _25601_ (.A1(_08427_),
    .A2(_06534_),
    .B1_N(_12189_),
    .X(_08428_));
 sky130_fd_sc_hd__clkbuf_8 _25602_ (.A(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__mux2_1 _25603_ (.A0(_07699_),
    .A1(net2227),
    .S(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__clkbuf_1 _25604_ (.A(_08430_),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_1 _25605_ (.A0(_07703_),
    .A1(net3116),
    .S(_08429_),
    .X(_08431_));
 sky130_fd_sc_hd__clkbuf_1 _25606_ (.A(_08431_),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _25607_ (.A0(_07705_),
    .A1(net2666),
    .S(_08429_),
    .X(_08432_));
 sky130_fd_sc_hd__clkbuf_1 _25608_ (.A(_08432_),
    .X(_02549_));
 sky130_fd_sc_hd__mux2_1 _25609_ (.A0(_07707_),
    .A1(net2459),
    .S(_08429_),
    .X(_08433_));
 sky130_fd_sc_hd__clkbuf_1 _25610_ (.A(_08433_),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _25611_ (.A0(_07709_),
    .A1(net3142),
    .S(_08429_),
    .X(_08434_));
 sky130_fd_sc_hd__clkbuf_1 _25612_ (.A(_08434_),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _25613_ (.A0(_07711_),
    .A1(net2786),
    .S(_08429_),
    .X(_08435_));
 sky130_fd_sc_hd__clkbuf_1 _25614_ (.A(_08435_),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _25615_ (.A0(_07713_),
    .A1(net2249),
    .S(_08429_),
    .X(_08436_));
 sky130_fd_sc_hd__clkbuf_1 _25616_ (.A(_08436_),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _25617_ (.A0(_07715_),
    .A1(net3490),
    .S(_08429_),
    .X(_08437_));
 sky130_fd_sc_hd__clkbuf_1 _25618_ (.A(_08437_),
    .X(_02554_));
 sky130_fd_sc_hd__buf_4 _25619_ (.A(_08427_),
    .X(_08438_));
 sky130_fd_sc_hd__buf_4 _25620_ (.A(_09125_),
    .X(_08439_));
 sky130_fd_sc_hd__buf_4 _25621_ (.A(_08427_),
    .X(_08440_));
 sky130_fd_sc_hd__nand2_1 _25622_ (.A(_08440_),
    .B(_12184_),
    .Y(_08441_));
 sky130_fd_sc_hd__o211a_1 _25623_ (.A1(_02850_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08441_),
    .X(_08442_));
 sky130_fd_sc_hd__mux2_1 _25624_ (.A0(_08442_),
    .A1(net2890),
    .S(_08429_),
    .X(_08443_));
 sky130_fd_sc_hd__clkbuf_1 _25625_ (.A(_08443_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _25626_ (.A(_08440_),
    .B(_12197_),
    .Y(_08444_));
 sky130_fd_sc_hd__o211a_1 _25627_ (.A1(_02860_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08444_),
    .X(_08445_));
 sky130_fd_sc_hd__mux2_1 _25628_ (.A0(_08445_),
    .A1(net2590),
    .S(_08429_),
    .X(_08446_));
 sky130_fd_sc_hd__clkbuf_1 _25629_ (.A(_08446_),
    .X(_02556_));
 sky130_fd_sc_hd__nand2_1 _25630_ (.A(_08440_),
    .B(_12205_),
    .Y(_08447_));
 sky130_fd_sc_hd__o211a_1 _25631_ (.A1(_02867_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08447_),
    .X(_08448_));
 sky130_fd_sc_hd__mux2_1 _25632_ (.A0(_08448_),
    .A1(net2983),
    .S(_08429_),
    .X(_08449_));
 sky130_fd_sc_hd__clkbuf_1 _25633_ (.A(_08449_),
    .X(_02557_));
 sky130_fd_sc_hd__nand2_1 _25634_ (.A(_08440_),
    .B(_12213_),
    .Y(_08450_));
 sky130_fd_sc_hd__o211a_1 _25635_ (.A1(_02874_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08450_),
    .X(_08451_));
 sky130_fd_sc_hd__mux2_1 _25636_ (.A0(_08451_),
    .A1(net2706),
    .S(_08429_),
    .X(_08452_));
 sky130_fd_sc_hd__clkbuf_1 _25637_ (.A(_08452_),
    .X(_02558_));
 sky130_fd_sc_hd__nand2_1 _25638_ (.A(_08440_),
    .B(_12221_),
    .Y(_08453_));
 sky130_fd_sc_hd__o211a_1 _25639_ (.A1(_02881_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__mux2_1 _25640_ (.A0(_08454_),
    .A1(net2757),
    .S(_08429_),
    .X(_08455_));
 sky130_fd_sc_hd__clkbuf_1 _25641_ (.A(_08455_),
    .X(_02559_));
 sky130_fd_sc_hd__nand2_1 _25642_ (.A(_08440_),
    .B(_12229_),
    .Y(_08456_));
 sky130_fd_sc_hd__o211a_1 _25643_ (.A1(_02888_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__mux2_1 _25644_ (.A0(_08457_),
    .A1(net2479),
    .S(_08429_),
    .X(_08458_));
 sky130_fd_sc_hd__clkbuf_1 _25645_ (.A(_08458_),
    .X(_02560_));
 sky130_fd_sc_hd__nand2_1 _25646_ (.A(_08440_),
    .B(_12237_),
    .Y(_08459_));
 sky130_fd_sc_hd__o211a_1 _25647_ (.A1(_02895_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__mux2_1 _25648_ (.A0(_08460_),
    .A1(net2646),
    .S(_08429_),
    .X(_08461_));
 sky130_fd_sc_hd__clkbuf_1 _25649_ (.A(_08461_),
    .X(_02561_));
 sky130_fd_sc_hd__nand2_1 _25650_ (.A(_08440_),
    .B(_12245_),
    .Y(_08462_));
 sky130_fd_sc_hd__o211a_1 _25651_ (.A1(_02902_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__mux2_1 _25652_ (.A0(_08463_),
    .A1(net3247),
    .S(_08429_),
    .X(_08464_));
 sky130_fd_sc_hd__clkbuf_1 _25653_ (.A(_08464_),
    .X(_02562_));
 sky130_fd_sc_hd__o211a_1 _25654_ (.A1(_02910_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08441_),
    .X(_08465_));
 sky130_fd_sc_hd__clkbuf_8 _25655_ (.A(_08428_),
    .X(_08466_));
 sky130_fd_sc_hd__mux2_1 _25656_ (.A0(_08465_),
    .A1(net3066),
    .S(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__clkbuf_1 _25657_ (.A(_08467_),
    .X(_02563_));
 sky130_fd_sc_hd__o211a_1 _25658_ (.A1(_02915_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08444_),
    .X(_08468_));
 sky130_fd_sc_hd__mux2_1 _25659_ (.A0(_08468_),
    .A1(net3354),
    .S(_08466_),
    .X(_08469_));
 sky130_fd_sc_hd__clkbuf_1 _25660_ (.A(_08469_),
    .X(_02564_));
 sky130_fd_sc_hd__o211a_1 _25661_ (.A1(_02920_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08447_),
    .X(_08470_));
 sky130_fd_sc_hd__mux2_1 _25662_ (.A0(_08470_),
    .A1(net3024),
    .S(_08466_),
    .X(_08471_));
 sky130_fd_sc_hd__clkbuf_1 _25663_ (.A(_08471_),
    .X(_02565_));
 sky130_fd_sc_hd__o211a_1 _25664_ (.A1(_02926_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08450_),
    .X(_08472_));
 sky130_fd_sc_hd__mux2_1 _25665_ (.A0(_08472_),
    .A1(net2330),
    .S(_08466_),
    .X(_08473_));
 sky130_fd_sc_hd__clkbuf_1 _25666_ (.A(_08473_),
    .X(_02566_));
 sky130_fd_sc_hd__o211a_1 _25667_ (.A1(_02931_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08453_),
    .X(_08474_));
 sky130_fd_sc_hd__mux2_1 _25668_ (.A0(_08474_),
    .A1(net3385),
    .S(_08466_),
    .X(_08475_));
 sky130_fd_sc_hd__clkbuf_1 _25669_ (.A(_08475_),
    .X(_02567_));
 sky130_fd_sc_hd__o211a_1 _25670_ (.A1(_02936_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08456_),
    .X(_08476_));
 sky130_fd_sc_hd__mux2_1 _25671_ (.A0(_08476_),
    .A1(net3154),
    .S(_08466_),
    .X(_08477_));
 sky130_fd_sc_hd__clkbuf_1 _25672_ (.A(_08477_),
    .X(_02568_));
 sky130_fd_sc_hd__o211a_1 _25673_ (.A1(_02941_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08459_),
    .X(_08478_));
 sky130_fd_sc_hd__mux2_1 _25674_ (.A0(_08478_),
    .A1(net2490),
    .S(_08466_),
    .X(_08479_));
 sky130_fd_sc_hd__clkbuf_1 _25675_ (.A(_08479_),
    .X(_02569_));
 sky130_fd_sc_hd__o211a_1 _25676_ (.A1(_02946_),
    .A2(_08438_),
    .B1(_08439_),
    .C1(_08462_),
    .X(_08480_));
 sky130_fd_sc_hd__mux2_1 _25677_ (.A0(_08480_),
    .A1(net2884),
    .S(_08466_),
    .X(_08481_));
 sky130_fd_sc_hd__clkbuf_1 _25678_ (.A(_08481_),
    .X(_02570_));
 sky130_fd_sc_hd__buf_4 _25679_ (.A(_09125_),
    .X(_08482_));
 sky130_fd_sc_hd__o211a_1 _25680_ (.A1(_12169_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08441_),
    .X(_08483_));
 sky130_fd_sc_hd__mux2_1 _25681_ (.A0(_08483_),
    .A1(net2681),
    .S(_08466_),
    .X(_08484_));
 sky130_fd_sc_hd__clkbuf_1 _25682_ (.A(_08484_),
    .X(_02571_));
 sky130_fd_sc_hd__o211a_1 _25683_ (.A1(_12194_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08444_),
    .X(_08485_));
 sky130_fd_sc_hd__mux2_1 _25684_ (.A0(_08485_),
    .A1(net3364),
    .S(_08466_),
    .X(_08486_));
 sky130_fd_sc_hd__clkbuf_1 _25685_ (.A(_08486_),
    .X(_02572_));
 sky130_fd_sc_hd__o211a_1 _25686_ (.A1(_12202_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08447_),
    .X(_08487_));
 sky130_fd_sc_hd__mux2_1 _25687_ (.A0(_08487_),
    .A1(net2527),
    .S(_08466_),
    .X(_08488_));
 sky130_fd_sc_hd__clkbuf_1 _25688_ (.A(_08488_),
    .X(_02573_));
 sky130_fd_sc_hd__o211a_1 _25689_ (.A1(_12210_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08450_),
    .X(_08489_));
 sky130_fd_sc_hd__mux2_1 _25690_ (.A0(_08489_),
    .A1(net2876),
    .S(_08466_),
    .X(_08490_));
 sky130_fd_sc_hd__clkbuf_1 _25691_ (.A(_08490_),
    .X(_02574_));
 sky130_fd_sc_hd__o211a_1 _25692_ (.A1(_12218_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08453_),
    .X(_08491_));
 sky130_fd_sc_hd__mux2_1 _25693_ (.A0(_08491_),
    .A1(net2422),
    .S(_08466_),
    .X(_08492_));
 sky130_fd_sc_hd__clkbuf_1 _25694_ (.A(_08492_),
    .X(_02575_));
 sky130_fd_sc_hd__o211a_1 _25695_ (.A1(_12226_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08456_),
    .X(_08493_));
 sky130_fd_sc_hd__mux2_1 _25696_ (.A0(_08493_),
    .A1(net2554),
    .S(_08466_),
    .X(_08494_));
 sky130_fd_sc_hd__clkbuf_1 _25697_ (.A(_08494_),
    .X(_02576_));
 sky130_fd_sc_hd__o211a_1 _25698_ (.A1(_12234_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08459_),
    .X(_08495_));
 sky130_fd_sc_hd__mux2_1 _25699_ (.A0(_08495_),
    .A1(net2360),
    .S(_08466_),
    .X(_08496_));
 sky130_fd_sc_hd__clkbuf_1 _25700_ (.A(_08496_),
    .X(_02577_));
 sky130_fd_sc_hd__o211a_1 _25701_ (.A1(_12242_),
    .A2(_08440_),
    .B1(_08482_),
    .C1(_08462_),
    .X(_08497_));
 sky130_fd_sc_hd__mux2_1 _25702_ (.A0(_08497_),
    .A1(net3160),
    .S(_08466_),
    .X(_08498_));
 sky130_fd_sc_hd__clkbuf_1 _25703_ (.A(_08498_),
    .X(_02578_));
 sky130_fd_sc_hd__nand2_1 _25704_ (.A(_03737_),
    .B(_12177_),
    .Y(_08499_));
 sky130_fd_sc_hd__a21bo_1 _25705_ (.A1(_08499_),
    .A2(_09109_),
    .B1_N(_12189_),
    .X(_08500_));
 sky130_fd_sc_hd__clkbuf_8 _25706_ (.A(_08500_),
    .X(_08501_));
 sky130_fd_sc_hd__mux2_1 _25707_ (.A0(_07699_),
    .A1(net3176),
    .S(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__clkbuf_1 _25708_ (.A(_08502_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _25709_ (.A0(_07703_),
    .A1(net3050),
    .S(_08501_),
    .X(_08503_));
 sky130_fd_sc_hd__clkbuf_1 _25710_ (.A(_08503_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _25711_ (.A0(_07705_),
    .A1(net3328),
    .S(_08501_),
    .X(_08504_));
 sky130_fd_sc_hd__clkbuf_1 _25712_ (.A(_08504_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _25713_ (.A0(_07707_),
    .A1(net2774),
    .S(_08501_),
    .X(_08505_));
 sky130_fd_sc_hd__clkbuf_1 _25714_ (.A(_08505_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _25715_ (.A0(_07709_),
    .A1(net2412),
    .S(_08501_),
    .X(_08506_));
 sky130_fd_sc_hd__clkbuf_1 _25716_ (.A(_08506_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _25717_ (.A0(_07711_),
    .A1(net2272),
    .S(_08501_),
    .X(_08507_));
 sky130_fd_sc_hd__clkbuf_1 _25718_ (.A(_08507_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _25719_ (.A0(_07713_),
    .A1(net3478),
    .S(_08501_),
    .X(_08508_));
 sky130_fd_sc_hd__clkbuf_1 _25720_ (.A(_08508_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _25721_ (.A0(_07715_),
    .A1(net3171),
    .S(_08501_),
    .X(_08509_));
 sky130_fd_sc_hd__clkbuf_1 _25722_ (.A(_08509_),
    .X(_02586_));
 sky130_fd_sc_hd__buf_4 _25723_ (.A(_08499_),
    .X(_08510_));
 sky130_fd_sc_hd__buf_4 _25724_ (.A(_08499_),
    .X(_08511_));
 sky130_fd_sc_hd__nand2_1 _25725_ (.A(_08511_),
    .B(_12184_),
    .Y(_08512_));
 sky130_fd_sc_hd__o211a_1 _25726_ (.A1(_02850_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08512_),
    .X(_08513_));
 sky130_fd_sc_hd__mux2_1 _25727_ (.A0(_08513_),
    .A1(net2308),
    .S(_08501_),
    .X(_08514_));
 sky130_fd_sc_hd__clkbuf_1 _25728_ (.A(_08514_),
    .X(_02587_));
 sky130_fd_sc_hd__nand2_1 _25729_ (.A(_08511_),
    .B(_12197_),
    .Y(_08515_));
 sky130_fd_sc_hd__o211a_1 _25730_ (.A1(_02860_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__mux2_1 _25731_ (.A0(_08516_),
    .A1(net3029),
    .S(_08501_),
    .X(_08517_));
 sky130_fd_sc_hd__clkbuf_1 _25732_ (.A(_08517_),
    .X(_02588_));
 sky130_fd_sc_hd__nand2_1 _25733_ (.A(_08511_),
    .B(_12205_),
    .Y(_08518_));
 sky130_fd_sc_hd__o211a_1 _25734_ (.A1(_02867_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__mux2_1 _25735_ (.A0(_08519_),
    .A1(net3167),
    .S(_08501_),
    .X(_08520_));
 sky130_fd_sc_hd__clkbuf_1 _25736_ (.A(_08520_),
    .X(_02589_));
 sky130_fd_sc_hd__nand2_1 _25737_ (.A(_08511_),
    .B(_12213_),
    .Y(_08521_));
 sky130_fd_sc_hd__o211a_1 _25738_ (.A1(_02874_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__mux2_1 _25739_ (.A0(_08522_),
    .A1(net2500),
    .S(_08501_),
    .X(_08523_));
 sky130_fd_sc_hd__clkbuf_1 _25740_ (.A(_08523_),
    .X(_02590_));
 sky130_fd_sc_hd__nand2_1 _25741_ (.A(_08511_),
    .B(_12221_),
    .Y(_08524_));
 sky130_fd_sc_hd__o211a_1 _25742_ (.A1(_02881_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__mux2_1 _25743_ (.A0(_08525_),
    .A1(net2678),
    .S(_08501_),
    .X(_08526_));
 sky130_fd_sc_hd__clkbuf_1 _25744_ (.A(_08526_),
    .X(_02591_));
 sky130_fd_sc_hd__nand2_1 _25745_ (.A(_08511_),
    .B(_12229_),
    .Y(_08527_));
 sky130_fd_sc_hd__o211a_1 _25746_ (.A1(_02888_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__mux2_1 _25747_ (.A0(_08528_),
    .A1(net2915),
    .S(_08501_),
    .X(_08529_));
 sky130_fd_sc_hd__clkbuf_1 _25748_ (.A(_08529_),
    .X(_02592_));
 sky130_fd_sc_hd__nand2_1 _25749_ (.A(_08511_),
    .B(_12237_),
    .Y(_08530_));
 sky130_fd_sc_hd__o211a_1 _25750_ (.A1(_02895_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__mux2_1 _25751_ (.A0(_08531_),
    .A1(net2728),
    .S(_08501_),
    .X(_08532_));
 sky130_fd_sc_hd__clkbuf_1 _25752_ (.A(_08532_),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_1 _25753_ (.A(_08511_),
    .B(_12245_),
    .Y(_08533_));
 sky130_fd_sc_hd__o211a_1 _25754_ (.A1(_02902_),
    .A2(_08510_),
    .B1(_08482_),
    .C1(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__mux2_1 _25755_ (.A0(_08534_),
    .A1(net3335),
    .S(_08501_),
    .X(_08535_));
 sky130_fd_sc_hd__clkbuf_1 _25756_ (.A(_08535_),
    .X(_02594_));
 sky130_fd_sc_hd__buf_4 _25757_ (.A(_09125_),
    .X(_08536_));
 sky130_fd_sc_hd__o211a_1 _25758_ (.A1(_02910_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08512_),
    .X(_08537_));
 sky130_fd_sc_hd__clkbuf_8 _25759_ (.A(_08500_),
    .X(_08538_));
 sky130_fd_sc_hd__mux2_1 _25760_ (.A0(_08537_),
    .A1(net2080),
    .S(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__clkbuf_1 _25761_ (.A(_08539_),
    .X(_02595_));
 sky130_fd_sc_hd__o211a_1 _25762_ (.A1(_02915_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08515_),
    .X(_08540_));
 sky130_fd_sc_hd__mux2_1 _25763_ (.A0(_08540_),
    .A1(net2079),
    .S(_08538_),
    .X(_08541_));
 sky130_fd_sc_hd__clkbuf_1 _25764_ (.A(_08541_),
    .X(_02596_));
 sky130_fd_sc_hd__o211a_1 _25765_ (.A1(_02920_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08518_),
    .X(_08542_));
 sky130_fd_sc_hd__mux2_1 _25766_ (.A0(_08542_),
    .A1(net2133),
    .S(_08538_),
    .X(_08543_));
 sky130_fd_sc_hd__clkbuf_1 _25767_ (.A(_08543_),
    .X(_02597_));
 sky130_fd_sc_hd__o211a_1 _25768_ (.A1(_02926_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08521_),
    .X(_08544_));
 sky130_fd_sc_hd__mux2_1 _25769_ (.A0(_08544_),
    .A1(net2452),
    .S(_08538_),
    .X(_08545_));
 sky130_fd_sc_hd__clkbuf_1 _25770_ (.A(_08545_),
    .X(_02598_));
 sky130_fd_sc_hd__o211a_1 _25771_ (.A1(_02931_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08524_),
    .X(_08546_));
 sky130_fd_sc_hd__mux2_1 _25772_ (.A0(_08546_),
    .A1(net2116),
    .S(_08538_),
    .X(_08547_));
 sky130_fd_sc_hd__clkbuf_1 _25773_ (.A(_08547_),
    .X(_02599_));
 sky130_fd_sc_hd__o211a_1 _25774_ (.A1(_02936_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08527_),
    .X(_08548_));
 sky130_fd_sc_hd__mux2_1 _25775_ (.A0(_08548_),
    .A1(net2091),
    .S(_08538_),
    .X(_08549_));
 sky130_fd_sc_hd__clkbuf_1 _25776_ (.A(_08549_),
    .X(_02600_));
 sky130_fd_sc_hd__o211a_1 _25777_ (.A1(_02941_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08530_),
    .X(_08550_));
 sky130_fd_sc_hd__mux2_1 _25778_ (.A0(_08550_),
    .A1(net2128),
    .S(_08538_),
    .X(_08551_));
 sky130_fd_sc_hd__clkbuf_1 _25779_ (.A(_08551_),
    .X(_02601_));
 sky130_fd_sc_hd__o211a_1 _25780_ (.A1(_02946_),
    .A2(_08510_),
    .B1(_08536_),
    .C1(_08533_),
    .X(_08552_));
 sky130_fd_sc_hd__mux2_1 _25781_ (.A0(_08552_),
    .A1(net2094),
    .S(_08538_),
    .X(_08553_));
 sky130_fd_sc_hd__clkbuf_1 _25782_ (.A(_08553_),
    .X(_02602_));
 sky130_fd_sc_hd__o211a_1 _25783_ (.A1(_12169_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08512_),
    .X(_08554_));
 sky130_fd_sc_hd__mux2_1 _25784_ (.A0(_08554_),
    .A1(net2698),
    .S(_08538_),
    .X(_08555_));
 sky130_fd_sc_hd__clkbuf_1 _25785_ (.A(_08555_),
    .X(_02603_));
 sky130_fd_sc_hd__o211a_1 _25786_ (.A1(_12194_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08515_),
    .X(_08556_));
 sky130_fd_sc_hd__mux2_1 _25787_ (.A0(_08556_),
    .A1(net3319),
    .S(_08538_),
    .X(_08557_));
 sky130_fd_sc_hd__clkbuf_1 _25788_ (.A(_08557_),
    .X(_02604_));
 sky130_fd_sc_hd__o211a_1 _25789_ (.A1(_12202_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08518_),
    .X(_08558_));
 sky130_fd_sc_hd__mux2_1 _25790_ (.A0(_08558_),
    .A1(net2578),
    .S(_08538_),
    .X(_08559_));
 sky130_fd_sc_hd__clkbuf_1 _25791_ (.A(_08559_),
    .X(_02605_));
 sky130_fd_sc_hd__o211a_1 _25792_ (.A1(_12210_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08521_),
    .X(_08560_));
 sky130_fd_sc_hd__mux2_1 _25793_ (.A0(_08560_),
    .A1(net2616),
    .S(_08538_),
    .X(_08561_));
 sky130_fd_sc_hd__clkbuf_1 _25794_ (.A(_08561_),
    .X(_02606_));
 sky130_fd_sc_hd__o211a_1 _25795_ (.A1(_12218_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08524_),
    .X(_08562_));
 sky130_fd_sc_hd__mux2_1 _25796_ (.A0(_08562_),
    .A1(net3211),
    .S(_08538_),
    .X(_08563_));
 sky130_fd_sc_hd__clkbuf_1 _25797_ (.A(_08563_),
    .X(_02607_));
 sky130_fd_sc_hd__o211a_1 _25798_ (.A1(_12226_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08527_),
    .X(_08564_));
 sky130_fd_sc_hd__mux2_1 _25799_ (.A0(_08564_),
    .A1(net2625),
    .S(_08538_),
    .X(_08565_));
 sky130_fd_sc_hd__clkbuf_1 _25800_ (.A(_08565_),
    .X(_02608_));
 sky130_fd_sc_hd__o211a_1 _25801_ (.A1(_12234_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08530_),
    .X(_08566_));
 sky130_fd_sc_hd__mux2_1 _25802_ (.A0(_08566_),
    .A1(net2597),
    .S(_08538_),
    .X(_08567_));
 sky130_fd_sc_hd__clkbuf_1 _25803_ (.A(_08567_),
    .X(_02609_));
 sky130_fd_sc_hd__o211a_1 _25804_ (.A1(_12242_),
    .A2(_08511_),
    .B1(_08536_),
    .C1(_08533_),
    .X(_08568_));
 sky130_fd_sc_hd__mux2_1 _25805_ (.A0(_08568_),
    .A1(net3071),
    .S(_08538_),
    .X(_08569_));
 sky130_fd_sc_hd__clkbuf_1 _25806_ (.A(_08569_),
    .X(_02610_));
 sky130_fd_sc_hd__nand2_1 _25807_ (.A(_03811_),
    .B(_12177_),
    .Y(_08570_));
 sky130_fd_sc_hd__a21bo_1 _25808_ (.A1(_08570_),
    .A2(_09109_),
    .B1_N(_12189_),
    .X(_08571_));
 sky130_fd_sc_hd__buf_6 _25809_ (.A(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__mux2_1 _25810_ (.A0(_07699_),
    .A1(net2385),
    .S(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__clkbuf_1 _25811_ (.A(_08573_),
    .X(_02611_));
 sky130_fd_sc_hd__mux2_1 _25812_ (.A0(_07703_),
    .A1(net3609),
    .S(_08572_),
    .X(_08574_));
 sky130_fd_sc_hd__clkbuf_1 _25813_ (.A(_08574_),
    .X(_02612_));
 sky130_fd_sc_hd__mux2_1 _25814_ (.A0(_07705_),
    .A1(net3533),
    .S(_08572_),
    .X(_08575_));
 sky130_fd_sc_hd__clkbuf_1 _25815_ (.A(_08575_),
    .X(_02613_));
 sky130_fd_sc_hd__mux2_1 _25816_ (.A0(_07707_),
    .A1(net2434),
    .S(_08572_),
    .X(_08576_));
 sky130_fd_sc_hd__clkbuf_1 _25817_ (.A(_08576_),
    .X(_02614_));
 sky130_fd_sc_hd__mux2_1 _25818_ (.A0(_07709_),
    .A1(net3222),
    .S(_08572_),
    .X(_08577_));
 sky130_fd_sc_hd__clkbuf_1 _25819_ (.A(_08577_),
    .X(_02615_));
 sky130_fd_sc_hd__mux2_1 _25820_ (.A0(_07711_),
    .A1(net3521),
    .S(_08572_),
    .X(_08578_));
 sky130_fd_sc_hd__clkbuf_1 _25821_ (.A(_08578_),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _25822_ (.A0(_07713_),
    .A1(net2321),
    .S(_08572_),
    .X(_08579_));
 sky130_fd_sc_hd__clkbuf_1 _25823_ (.A(_08579_),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_1 _25824_ (.A0(_07715_),
    .A1(net2626),
    .S(_08572_),
    .X(_08580_));
 sky130_fd_sc_hd__clkbuf_1 _25825_ (.A(_08580_),
    .X(_02618_));
 sky130_fd_sc_hd__buf_4 _25826_ (.A(_08570_),
    .X(_08581_));
 sky130_fd_sc_hd__buf_4 _25827_ (.A(_09125_),
    .X(_08582_));
 sky130_fd_sc_hd__buf_4 _25828_ (.A(_08570_),
    .X(_08583_));
 sky130_fd_sc_hd__nand2_1 _25829_ (.A(_08583_),
    .B(_12184_),
    .Y(_08584_));
 sky130_fd_sc_hd__o211a_1 _25830_ (.A1(_02850_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__mux2_1 _25831_ (.A0(_08585_),
    .A1(net3776),
    .S(_08572_),
    .X(_08586_));
 sky130_fd_sc_hd__clkbuf_1 _25832_ (.A(_08586_),
    .X(_02619_));
 sky130_fd_sc_hd__nand2_1 _25833_ (.A(_08583_),
    .B(_12197_),
    .Y(_08587_));
 sky130_fd_sc_hd__o211a_1 _25834_ (.A1(_02860_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08587_),
    .X(_08588_));
 sky130_fd_sc_hd__mux2_1 _25835_ (.A0(_08588_),
    .A1(net2240),
    .S(_08572_),
    .X(_08589_));
 sky130_fd_sc_hd__clkbuf_1 _25836_ (.A(_08589_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_1 _25837_ (.A(_08583_),
    .B(_12205_),
    .Y(_08590_));
 sky130_fd_sc_hd__o211a_1 _25838_ (.A1(_02867_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__mux2_1 _25839_ (.A0(_08591_),
    .A1(net3384),
    .S(_08572_),
    .X(_08592_));
 sky130_fd_sc_hd__clkbuf_1 _25840_ (.A(_08592_),
    .X(_02621_));
 sky130_fd_sc_hd__nand2_1 _25841_ (.A(_08583_),
    .B(_12213_),
    .Y(_08593_));
 sky130_fd_sc_hd__o211a_1 _25842_ (.A1(_02874_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08593_),
    .X(_08594_));
 sky130_fd_sc_hd__mux2_1 _25843_ (.A0(_08594_),
    .A1(net3111),
    .S(_08572_),
    .X(_08595_));
 sky130_fd_sc_hd__clkbuf_1 _25844_ (.A(_08595_),
    .X(_02622_));
 sky130_fd_sc_hd__nand2_1 _25845_ (.A(_08583_),
    .B(_12221_),
    .Y(_08596_));
 sky130_fd_sc_hd__o211a_1 _25846_ (.A1(_02881_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__mux2_1 _25847_ (.A0(_08597_),
    .A1(net2487),
    .S(_08572_),
    .X(_08598_));
 sky130_fd_sc_hd__clkbuf_1 _25848_ (.A(_08598_),
    .X(_02623_));
 sky130_fd_sc_hd__nand2_1 _25849_ (.A(_08583_),
    .B(_12229_),
    .Y(_08599_));
 sky130_fd_sc_hd__o211a_1 _25850_ (.A1(_02888_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__mux2_1 _25851_ (.A0(_08600_),
    .A1(net3094),
    .S(_08572_),
    .X(_08601_));
 sky130_fd_sc_hd__clkbuf_1 _25852_ (.A(_08601_),
    .X(_02624_));
 sky130_fd_sc_hd__nand2_1 _25853_ (.A(_08583_),
    .B(_12237_),
    .Y(_08602_));
 sky130_fd_sc_hd__o211a_1 _25854_ (.A1(_02895_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__mux2_1 _25855_ (.A0(_08603_),
    .A1(net3655),
    .S(_08572_),
    .X(_08604_));
 sky130_fd_sc_hd__clkbuf_1 _25856_ (.A(_08604_),
    .X(_02625_));
 sky130_fd_sc_hd__nand2_1 _25857_ (.A(_08583_),
    .B(_12245_),
    .Y(_08605_));
 sky130_fd_sc_hd__o211a_1 _25858_ (.A1(_02902_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__mux2_1 _25859_ (.A0(_08606_),
    .A1(net3761),
    .S(_08572_),
    .X(_08607_));
 sky130_fd_sc_hd__clkbuf_1 _25860_ (.A(_08607_),
    .X(_02626_));
 sky130_fd_sc_hd__o211a_1 _25861_ (.A1(_02910_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08584_),
    .X(_08608_));
 sky130_fd_sc_hd__clkbuf_8 _25862_ (.A(_08571_),
    .X(_08609_));
 sky130_fd_sc_hd__mux2_1 _25863_ (.A0(_08608_),
    .A1(net2518),
    .S(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__clkbuf_1 _25864_ (.A(_08610_),
    .X(_02627_));
 sky130_fd_sc_hd__o211a_1 _25865_ (.A1(_02915_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08587_),
    .X(_08611_));
 sky130_fd_sc_hd__mux2_1 _25866_ (.A0(_08611_),
    .A1(net2758),
    .S(_08609_),
    .X(_08612_));
 sky130_fd_sc_hd__clkbuf_1 _25867_ (.A(_08612_),
    .X(_02628_));
 sky130_fd_sc_hd__o211a_1 _25868_ (.A1(_02920_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08590_),
    .X(_08613_));
 sky130_fd_sc_hd__mux2_1 _25869_ (.A0(_08613_),
    .A1(net3074),
    .S(_08609_),
    .X(_08614_));
 sky130_fd_sc_hd__clkbuf_1 _25870_ (.A(_08614_),
    .X(_02629_));
 sky130_fd_sc_hd__o211a_1 _25871_ (.A1(_02926_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08593_),
    .X(_08615_));
 sky130_fd_sc_hd__mux2_1 _25872_ (.A0(_08615_),
    .A1(net2544),
    .S(_08609_),
    .X(_08616_));
 sky130_fd_sc_hd__clkbuf_1 _25873_ (.A(_08616_),
    .X(_02630_));
 sky130_fd_sc_hd__o211a_1 _25874_ (.A1(_02931_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08596_),
    .X(_08617_));
 sky130_fd_sc_hd__mux2_1 _25875_ (.A0(_08617_),
    .A1(net3240),
    .S(_08609_),
    .X(_08618_));
 sky130_fd_sc_hd__clkbuf_1 _25876_ (.A(_08618_),
    .X(_02631_));
 sky130_fd_sc_hd__o211a_1 _25877_ (.A1(_02936_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08599_),
    .X(_08619_));
 sky130_fd_sc_hd__mux2_1 _25878_ (.A0(_08619_),
    .A1(net2821),
    .S(_08609_),
    .X(_08620_));
 sky130_fd_sc_hd__clkbuf_1 _25879_ (.A(_08620_),
    .X(_02632_));
 sky130_fd_sc_hd__o211a_1 _25880_ (.A1(_02941_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08602_),
    .X(_08621_));
 sky130_fd_sc_hd__mux2_1 _25881_ (.A0(_08621_),
    .A1(net3286),
    .S(_08609_),
    .X(_08622_));
 sky130_fd_sc_hd__clkbuf_1 _25882_ (.A(_08622_),
    .X(_02633_));
 sky130_fd_sc_hd__o211a_1 _25883_ (.A1(_02946_),
    .A2(_08581_),
    .B1(_08582_),
    .C1(_08605_),
    .X(_08623_));
 sky130_fd_sc_hd__mux2_1 _25884_ (.A0(_08623_),
    .A1(net3281),
    .S(_08609_),
    .X(_08624_));
 sky130_fd_sc_hd__clkbuf_1 _25885_ (.A(_08624_),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_8 _25886_ (.A(_09125_),
    .X(_08625_));
 sky130_fd_sc_hd__o211a_1 _25887_ (.A1(_12169_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08584_),
    .X(_08626_));
 sky130_fd_sc_hd__mux2_1 _25888_ (.A0(_08626_),
    .A1(net2954),
    .S(_08609_),
    .X(_08627_));
 sky130_fd_sc_hd__clkbuf_1 _25889_ (.A(_08627_),
    .X(_02635_));
 sky130_fd_sc_hd__o211a_1 _25890_ (.A1(_12194_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08587_),
    .X(_08628_));
 sky130_fd_sc_hd__mux2_1 _25891_ (.A0(_08628_),
    .A1(net2541),
    .S(_08609_),
    .X(_08629_));
 sky130_fd_sc_hd__clkbuf_1 _25892_ (.A(_08629_),
    .X(_02636_));
 sky130_fd_sc_hd__o211a_1 _25893_ (.A1(_12202_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08590_),
    .X(_08630_));
 sky130_fd_sc_hd__mux2_1 _25894_ (.A0(_08630_),
    .A1(net2135),
    .S(_08609_),
    .X(_08631_));
 sky130_fd_sc_hd__clkbuf_1 _25895_ (.A(_08631_),
    .X(_02637_));
 sky130_fd_sc_hd__o211a_1 _25896_ (.A1(_12210_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08593_),
    .X(_08632_));
 sky130_fd_sc_hd__mux2_1 _25897_ (.A0(_08632_),
    .A1(net2569),
    .S(_08609_),
    .X(_08633_));
 sky130_fd_sc_hd__clkbuf_1 _25898_ (.A(_08633_),
    .X(_02638_));
 sky130_fd_sc_hd__o211a_1 _25899_ (.A1(_12218_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08596_),
    .X(_08634_));
 sky130_fd_sc_hd__mux2_1 _25900_ (.A0(_08634_),
    .A1(net2644),
    .S(_08609_),
    .X(_08635_));
 sky130_fd_sc_hd__clkbuf_1 _25901_ (.A(_08635_),
    .X(_02639_));
 sky130_fd_sc_hd__o211a_1 _25902_ (.A1(_12226_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08599_),
    .X(_08636_));
 sky130_fd_sc_hd__mux2_1 _25903_ (.A0(_08636_),
    .A1(net2694),
    .S(_08609_),
    .X(_08637_));
 sky130_fd_sc_hd__clkbuf_1 _25904_ (.A(_08637_),
    .X(_02640_));
 sky130_fd_sc_hd__o211a_1 _25905_ (.A1(_12234_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08602_),
    .X(_08638_));
 sky130_fd_sc_hd__mux2_1 _25906_ (.A0(_08638_),
    .A1(net2892),
    .S(_08609_),
    .X(_08639_));
 sky130_fd_sc_hd__clkbuf_1 _25907_ (.A(_08639_),
    .X(_02641_));
 sky130_fd_sc_hd__o211a_1 _25908_ (.A1(_12242_),
    .A2(_08583_),
    .B1(_08625_),
    .C1(_08605_),
    .X(_08640_));
 sky130_fd_sc_hd__mux2_1 _25909_ (.A0(_08640_),
    .A1(net2571),
    .S(_08609_),
    .X(_08641_));
 sky130_fd_sc_hd__clkbuf_1 _25910_ (.A(_08641_),
    .X(_02642_));
 sky130_fd_sc_hd__nand2_1 _25911_ (.A(_03884_),
    .B(_12177_),
    .Y(_08642_));
 sky130_fd_sc_hd__a21bo_1 _25912_ (.A1(_08642_),
    .A2(_09109_),
    .B1_N(_12189_),
    .X(_08643_));
 sky130_fd_sc_hd__clkbuf_8 _25913_ (.A(_08643_),
    .X(_08644_));
 sky130_fd_sc_hd__mux2_1 _25914_ (.A0(_07699_),
    .A1(net2320),
    .S(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__clkbuf_1 _25915_ (.A(_08645_),
    .X(_02643_));
 sky130_fd_sc_hd__mux2_1 _25916_ (.A0(_07703_),
    .A1(net3392),
    .S(_08644_),
    .X(_08646_));
 sky130_fd_sc_hd__clkbuf_1 _25917_ (.A(_08646_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _25918_ (.A0(_07705_),
    .A1(net2618),
    .S(_08644_),
    .X(_08647_));
 sky130_fd_sc_hd__clkbuf_1 _25919_ (.A(_08647_),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _25920_ (.A0(_07707_),
    .A1(net2791),
    .S(_08644_),
    .X(_08648_));
 sky130_fd_sc_hd__clkbuf_1 _25921_ (.A(_08648_),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _25922_ (.A0(_07709_),
    .A1(net2832),
    .S(_08644_),
    .X(_08649_));
 sky130_fd_sc_hd__clkbuf_1 _25923_ (.A(_08649_),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _25924_ (.A0(_07711_),
    .A1(net2718),
    .S(_08644_),
    .X(_08650_));
 sky130_fd_sc_hd__clkbuf_1 _25925_ (.A(_08650_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_1 _25926_ (.A0(_07713_),
    .A1(net3232),
    .S(_08644_),
    .X(_08651_));
 sky130_fd_sc_hd__clkbuf_1 _25927_ (.A(_08651_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _25928_ (.A0(_07715_),
    .A1(net2261),
    .S(_08644_),
    .X(_08652_));
 sky130_fd_sc_hd__clkbuf_1 _25929_ (.A(_08652_),
    .X(_02650_));
 sky130_fd_sc_hd__buf_4 _25930_ (.A(_08642_),
    .X(_08653_));
 sky130_fd_sc_hd__buf_4 _25931_ (.A(_08642_),
    .X(_08654_));
 sky130_fd_sc_hd__nand2_1 _25932_ (.A(_08654_),
    .B(_12184_),
    .Y(_08655_));
 sky130_fd_sc_hd__o211a_1 _25933_ (.A1(_02850_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08655_),
    .X(_08656_));
 sky130_fd_sc_hd__mux2_1 _25934_ (.A0(_08656_),
    .A1(net2624),
    .S(_08644_),
    .X(_08657_));
 sky130_fd_sc_hd__clkbuf_1 _25935_ (.A(_08657_),
    .X(_02651_));
 sky130_fd_sc_hd__nand2_1 _25936_ (.A(_08654_),
    .B(_12197_),
    .Y(_08658_));
 sky130_fd_sc_hd__o211a_1 _25937_ (.A1(_02860_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08658_),
    .X(_08659_));
 sky130_fd_sc_hd__mux2_1 _25938_ (.A0(_08659_),
    .A1(net2572),
    .S(_08644_),
    .X(_08660_));
 sky130_fd_sc_hd__clkbuf_1 _25939_ (.A(_08660_),
    .X(_02652_));
 sky130_fd_sc_hd__nand2_1 _25940_ (.A(_08654_),
    .B(_12205_),
    .Y(_08661_));
 sky130_fd_sc_hd__o211a_1 _25941_ (.A1(_02867_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08661_),
    .X(_08662_));
 sky130_fd_sc_hd__mux2_1 _25942_ (.A0(_08662_),
    .A1(net3576),
    .S(_08644_),
    .X(_08663_));
 sky130_fd_sc_hd__clkbuf_1 _25943_ (.A(_08663_),
    .X(_02653_));
 sky130_fd_sc_hd__nand2_1 _25944_ (.A(_08654_),
    .B(_12213_),
    .Y(_08664_));
 sky130_fd_sc_hd__o211a_1 _25945_ (.A1(_02874_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08664_),
    .X(_08665_));
 sky130_fd_sc_hd__mux2_1 _25946_ (.A0(_08665_),
    .A1(net3429),
    .S(_08644_),
    .X(_08666_));
 sky130_fd_sc_hd__clkbuf_1 _25947_ (.A(_08666_),
    .X(_02654_));
 sky130_fd_sc_hd__nand2_1 _25948_ (.A(_08654_),
    .B(_12221_),
    .Y(_08667_));
 sky130_fd_sc_hd__o211a_1 _25949_ (.A1(_02881_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08667_),
    .X(_08668_));
 sky130_fd_sc_hd__mux2_1 _25950_ (.A0(_08668_),
    .A1(net2424),
    .S(_08644_),
    .X(_08669_));
 sky130_fd_sc_hd__clkbuf_1 _25951_ (.A(_08669_),
    .X(_02655_));
 sky130_fd_sc_hd__nand2_1 _25952_ (.A(_08654_),
    .B(_12229_),
    .Y(_08670_));
 sky130_fd_sc_hd__o211a_1 _25953_ (.A1(_02888_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08670_),
    .X(_08671_));
 sky130_fd_sc_hd__mux2_1 _25954_ (.A0(_08671_),
    .A1(net2373),
    .S(_08644_),
    .X(_08672_));
 sky130_fd_sc_hd__clkbuf_1 _25955_ (.A(_08672_),
    .X(_02656_));
 sky130_fd_sc_hd__nand2_1 _25956_ (.A(_08654_),
    .B(_12237_),
    .Y(_08673_));
 sky130_fd_sc_hd__o211a_1 _25957_ (.A1(_02895_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08673_),
    .X(_08674_));
 sky130_fd_sc_hd__mux2_1 _25958_ (.A0(_08674_),
    .A1(net2938),
    .S(_08644_),
    .X(_08675_));
 sky130_fd_sc_hd__clkbuf_1 _25959_ (.A(_08675_),
    .X(_02657_));
 sky130_fd_sc_hd__nand2_1 _25960_ (.A(_08654_),
    .B(_12245_),
    .Y(_08676_));
 sky130_fd_sc_hd__o211a_1 _25961_ (.A1(_02902_),
    .A2(_08653_),
    .B1(_08625_),
    .C1(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__mux2_1 _25962_ (.A0(_08677_),
    .A1(net3195),
    .S(_08644_),
    .X(_08678_));
 sky130_fd_sc_hd__clkbuf_1 _25963_ (.A(_08678_),
    .X(_02658_));
 sky130_fd_sc_hd__buf_4 _25964_ (.A(_09125_),
    .X(_08679_));
 sky130_fd_sc_hd__o211a_1 _25965_ (.A1(_02910_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08655_),
    .X(_08680_));
 sky130_fd_sc_hd__clkbuf_8 _25966_ (.A(_08643_),
    .X(_08681_));
 sky130_fd_sc_hd__mux2_1 _25967_ (.A0(_08680_),
    .A1(net2927),
    .S(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__clkbuf_1 _25968_ (.A(_08682_),
    .X(_02659_));
 sky130_fd_sc_hd__o211a_1 _25969_ (.A1(_02915_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08658_),
    .X(_08683_));
 sky130_fd_sc_hd__mux2_1 _25970_ (.A0(_08683_),
    .A1(net2558),
    .S(_08681_),
    .X(_08684_));
 sky130_fd_sc_hd__clkbuf_1 _25971_ (.A(_08684_),
    .X(_02660_));
 sky130_fd_sc_hd__o211a_1 _25972_ (.A1(_02920_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08661_),
    .X(_08685_));
 sky130_fd_sc_hd__mux2_1 _25973_ (.A0(_08685_),
    .A1(net2994),
    .S(_08681_),
    .X(_08686_));
 sky130_fd_sc_hd__clkbuf_1 _25974_ (.A(_08686_),
    .X(_02661_));
 sky130_fd_sc_hd__o211a_1 _25975_ (.A1(_02926_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08664_),
    .X(_08687_));
 sky130_fd_sc_hd__mux2_1 _25976_ (.A0(_08687_),
    .A1(net2878),
    .S(_08681_),
    .X(_08688_));
 sky130_fd_sc_hd__clkbuf_1 _25977_ (.A(_08688_),
    .X(_02662_));
 sky130_fd_sc_hd__o211a_1 _25978_ (.A1(_02931_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08667_),
    .X(_08689_));
 sky130_fd_sc_hd__mux2_1 _25979_ (.A0(_08689_),
    .A1(net2469),
    .S(_08681_),
    .X(_08690_));
 sky130_fd_sc_hd__clkbuf_1 _25980_ (.A(_08690_),
    .X(_02663_));
 sky130_fd_sc_hd__o211a_1 _25981_ (.A1(_02936_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08670_),
    .X(_08691_));
 sky130_fd_sc_hd__mux2_1 _25982_ (.A0(_08691_),
    .A1(net3133),
    .S(_08681_),
    .X(_08692_));
 sky130_fd_sc_hd__clkbuf_1 _25983_ (.A(_08692_),
    .X(_02664_));
 sky130_fd_sc_hd__o211a_1 _25984_ (.A1(_02941_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08673_),
    .X(_08693_));
 sky130_fd_sc_hd__mux2_1 _25985_ (.A0(_08693_),
    .A1(net3251),
    .S(_08681_),
    .X(_08694_));
 sky130_fd_sc_hd__clkbuf_1 _25986_ (.A(_08694_),
    .X(_02665_));
 sky130_fd_sc_hd__o211a_1 _25987_ (.A1(_02946_),
    .A2(_08653_),
    .B1(_08679_),
    .C1(_08676_),
    .X(_08695_));
 sky130_fd_sc_hd__mux2_1 _25988_ (.A0(_08695_),
    .A1(net2827),
    .S(_08681_),
    .X(_08696_));
 sky130_fd_sc_hd__clkbuf_1 _25989_ (.A(_08696_),
    .X(_02666_));
 sky130_fd_sc_hd__o211a_1 _25990_ (.A1(_12169_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08655_),
    .X(_08697_));
 sky130_fd_sc_hd__mux2_1 _25991_ (.A0(_08697_),
    .A1(net3372),
    .S(_08681_),
    .X(_08698_));
 sky130_fd_sc_hd__clkbuf_1 _25992_ (.A(_08698_),
    .X(_02667_));
 sky130_fd_sc_hd__o211a_1 _25993_ (.A1(_12194_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08658_),
    .X(_08699_));
 sky130_fd_sc_hd__mux2_1 _25994_ (.A0(_08699_),
    .A1(net2386),
    .S(_08681_),
    .X(_08700_));
 sky130_fd_sc_hd__clkbuf_1 _25995_ (.A(_08700_),
    .X(_02668_));
 sky130_fd_sc_hd__o211a_1 _25996_ (.A1(_12202_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08661_),
    .X(_08701_));
 sky130_fd_sc_hd__mux2_1 _25997_ (.A0(_08701_),
    .A1(net2730),
    .S(_08681_),
    .X(_08702_));
 sky130_fd_sc_hd__clkbuf_1 _25998_ (.A(_08702_),
    .X(_02669_));
 sky130_fd_sc_hd__o211a_1 _25999_ (.A1(_12210_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08664_),
    .X(_08703_));
 sky130_fd_sc_hd__mux2_1 _26000_ (.A0(_08703_),
    .A1(net2623),
    .S(_08681_),
    .X(_08704_));
 sky130_fd_sc_hd__clkbuf_1 _26001_ (.A(_08704_),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_1 _26002_ (.A1(_12218_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08667_),
    .X(_08705_));
 sky130_fd_sc_hd__mux2_1 _26003_ (.A0(_08705_),
    .A1(net3047),
    .S(_08681_),
    .X(_08706_));
 sky130_fd_sc_hd__clkbuf_1 _26004_ (.A(_08706_),
    .X(_02671_));
 sky130_fd_sc_hd__o211a_1 _26005_ (.A1(_12226_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08670_),
    .X(_08707_));
 sky130_fd_sc_hd__mux2_1 _26006_ (.A0(_08707_),
    .A1(net3059),
    .S(_08681_),
    .X(_08708_));
 sky130_fd_sc_hd__clkbuf_1 _26007_ (.A(_08708_),
    .X(_02672_));
 sky130_fd_sc_hd__o211a_1 _26008_ (.A1(_12234_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08673_),
    .X(_08709_));
 sky130_fd_sc_hd__mux2_1 _26009_ (.A0(_08709_),
    .A1(net2709),
    .S(_08681_),
    .X(_08710_));
 sky130_fd_sc_hd__clkbuf_1 _26010_ (.A(_08710_),
    .X(_02673_));
 sky130_fd_sc_hd__o211a_1 _26011_ (.A1(_12242_),
    .A2(_08654_),
    .B1(_08679_),
    .C1(_08676_),
    .X(_08711_));
 sky130_fd_sc_hd__mux2_1 _26012_ (.A0(_08711_),
    .A1(net2974),
    .S(_08681_),
    .X(_08712_));
 sky130_fd_sc_hd__clkbuf_1 _26013_ (.A(_08712_),
    .X(_02674_));
 sky130_fd_sc_hd__nand2_1 _26014_ (.A(_03957_),
    .B(_12177_),
    .Y(_08713_));
 sky130_fd_sc_hd__a21bo_1 _26015_ (.A1(_08713_),
    .A2(_09109_),
    .B1_N(_12189_),
    .X(_08714_));
 sky130_fd_sc_hd__buf_6 _26016_ (.A(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__mux2_1 _26017_ (.A0(_07699_),
    .A1(net3530),
    .S(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__clkbuf_1 _26018_ (.A(_08716_),
    .X(_02675_));
 sky130_fd_sc_hd__mux2_1 _26019_ (.A0(_07703_),
    .A1(net3479),
    .S(_08715_),
    .X(_08717_));
 sky130_fd_sc_hd__clkbuf_1 _26020_ (.A(_08717_),
    .X(_02676_));
 sky130_fd_sc_hd__mux2_1 _26021_ (.A0(_07705_),
    .A1(net3022),
    .S(_08715_),
    .X(_08718_));
 sky130_fd_sc_hd__clkbuf_1 _26022_ (.A(_08718_),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _26023_ (.A0(_07707_),
    .A1(net2450),
    .S(_08715_),
    .X(_08719_));
 sky130_fd_sc_hd__clkbuf_1 _26024_ (.A(_08719_),
    .X(_02678_));
 sky130_fd_sc_hd__mux2_1 _26025_ (.A0(_07709_),
    .A1(net2484),
    .S(_08715_),
    .X(_08720_));
 sky130_fd_sc_hd__clkbuf_1 _26026_ (.A(_08720_),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _26027_ (.A0(_07711_),
    .A1(net3237),
    .S(_08715_),
    .X(_08721_));
 sky130_fd_sc_hd__clkbuf_1 _26028_ (.A(_08721_),
    .X(_02680_));
 sky130_fd_sc_hd__mux2_1 _26029_ (.A0(_07713_),
    .A1(net3468),
    .S(_08715_),
    .X(_08722_));
 sky130_fd_sc_hd__clkbuf_1 _26030_ (.A(_08722_),
    .X(_02681_));
 sky130_fd_sc_hd__mux2_1 _26031_ (.A0(_07715_),
    .A1(net2224),
    .S(_08715_),
    .X(_08723_));
 sky130_fd_sc_hd__clkbuf_1 _26032_ (.A(_08723_),
    .X(_02682_));
 sky130_fd_sc_hd__buf_4 _26033_ (.A(_08713_),
    .X(_08724_));
 sky130_fd_sc_hd__buf_4 _26034_ (.A(_09125_),
    .X(_08725_));
 sky130_fd_sc_hd__buf_4 _26035_ (.A(_08713_),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_1 _26036_ (.A(_08726_),
    .B(_12184_),
    .Y(_08727_));
 sky130_fd_sc_hd__o211a_1 _26037_ (.A1(_02850_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08727_),
    .X(_08728_));
 sky130_fd_sc_hd__mux2_1 _26038_ (.A0(_08728_),
    .A1(net3037),
    .S(_08715_),
    .X(_08729_));
 sky130_fd_sc_hd__clkbuf_1 _26039_ (.A(_08729_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _26040_ (.A(_08726_),
    .B(_12197_),
    .Y(_08730_));
 sky130_fd_sc_hd__o211a_1 _26041_ (.A1(_02860_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08730_),
    .X(_08731_));
 sky130_fd_sc_hd__mux2_1 _26042_ (.A0(_08731_),
    .A1(net2150),
    .S(_08715_),
    .X(_08732_));
 sky130_fd_sc_hd__clkbuf_1 _26043_ (.A(_08732_),
    .X(_02684_));
 sky130_fd_sc_hd__nand2_1 _26044_ (.A(_08726_),
    .B(_12205_),
    .Y(_08733_));
 sky130_fd_sc_hd__o211a_1 _26045_ (.A1(_02867_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__mux2_1 _26046_ (.A0(_08734_),
    .A1(net2740),
    .S(_08715_),
    .X(_08735_));
 sky130_fd_sc_hd__clkbuf_1 _26047_ (.A(_08735_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_1 _26048_ (.A(_08726_),
    .B(_12213_),
    .Y(_08736_));
 sky130_fd_sc_hd__o211a_1 _26049_ (.A1(_02874_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08736_),
    .X(_08737_));
 sky130_fd_sc_hd__mux2_1 _26050_ (.A0(_08737_),
    .A1(net2534),
    .S(_08715_),
    .X(_08738_));
 sky130_fd_sc_hd__clkbuf_1 _26051_ (.A(_08738_),
    .X(_02686_));
 sky130_fd_sc_hd__nand2_1 _26052_ (.A(_08726_),
    .B(_12221_),
    .Y(_08739_));
 sky130_fd_sc_hd__o211a_1 _26053_ (.A1(_02881_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08739_),
    .X(_08740_));
 sky130_fd_sc_hd__mux2_1 _26054_ (.A0(_08740_),
    .A1(net2280),
    .S(_08715_),
    .X(_08741_));
 sky130_fd_sc_hd__clkbuf_1 _26055_ (.A(_08741_),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_1 _26056_ (.A(_08726_),
    .B(_12229_),
    .Y(_08742_));
 sky130_fd_sc_hd__o211a_1 _26057_ (.A1(_02888_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__mux2_1 _26058_ (.A0(_08743_),
    .A1(net3303),
    .S(_08715_),
    .X(_08744_));
 sky130_fd_sc_hd__clkbuf_1 _26059_ (.A(_08744_),
    .X(_02688_));
 sky130_fd_sc_hd__nand2_1 _26060_ (.A(_08726_),
    .B(_12237_),
    .Y(_08745_));
 sky130_fd_sc_hd__o211a_1 _26061_ (.A1(_02895_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08745_),
    .X(_08746_));
 sky130_fd_sc_hd__mux2_1 _26062_ (.A0(_08746_),
    .A1(net2766),
    .S(_08715_),
    .X(_08747_));
 sky130_fd_sc_hd__clkbuf_1 _26063_ (.A(_08747_),
    .X(_02689_));
 sky130_fd_sc_hd__nand2_1 _26064_ (.A(_08726_),
    .B(_12245_),
    .Y(_08748_));
 sky130_fd_sc_hd__o211a_1 _26065_ (.A1(_02902_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__mux2_1 _26066_ (.A0(_08749_),
    .A1(net2517),
    .S(_08715_),
    .X(_08750_));
 sky130_fd_sc_hd__clkbuf_1 _26067_ (.A(_08750_),
    .X(_02690_));
 sky130_fd_sc_hd__o211a_1 _26068_ (.A1(_02910_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08727_),
    .X(_08751_));
 sky130_fd_sc_hd__clkbuf_8 _26069_ (.A(_08714_),
    .X(_08752_));
 sky130_fd_sc_hd__mux2_1 _26070_ (.A0(_08751_),
    .A1(net3005),
    .S(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__clkbuf_1 _26071_ (.A(_08753_),
    .X(_02691_));
 sky130_fd_sc_hd__o211a_1 _26072_ (.A1(_02915_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08730_),
    .X(_08754_));
 sky130_fd_sc_hd__mux2_1 _26073_ (.A0(_08754_),
    .A1(net2390),
    .S(_08752_),
    .X(_08755_));
 sky130_fd_sc_hd__clkbuf_1 _26074_ (.A(_08755_),
    .X(_02692_));
 sky130_fd_sc_hd__o211a_1 _26075_ (.A1(_02920_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08733_),
    .X(_08756_));
 sky130_fd_sc_hd__mux2_1 _26076_ (.A0(_08756_),
    .A1(net3326),
    .S(_08752_),
    .X(_08757_));
 sky130_fd_sc_hd__clkbuf_1 _26077_ (.A(_08757_),
    .X(_02693_));
 sky130_fd_sc_hd__o211a_1 _26078_ (.A1(_02926_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08736_),
    .X(_08758_));
 sky130_fd_sc_hd__mux2_1 _26079_ (.A0(_08758_),
    .A1(net2598),
    .S(_08752_),
    .X(_08759_));
 sky130_fd_sc_hd__clkbuf_1 _26080_ (.A(_08759_),
    .X(_02694_));
 sky130_fd_sc_hd__o211a_1 _26081_ (.A1(_02931_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08739_),
    .X(_08760_));
 sky130_fd_sc_hd__mux2_1 _26082_ (.A0(_08760_),
    .A1(net2660),
    .S(_08752_),
    .X(_08761_));
 sky130_fd_sc_hd__clkbuf_1 _26083_ (.A(_08761_),
    .X(_02695_));
 sky130_fd_sc_hd__o211a_1 _26084_ (.A1(_02936_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08742_),
    .X(_08762_));
 sky130_fd_sc_hd__mux2_1 _26085_ (.A0(_08762_),
    .A1(net2667),
    .S(_08752_),
    .X(_08763_));
 sky130_fd_sc_hd__clkbuf_1 _26086_ (.A(_08763_),
    .X(_02696_));
 sky130_fd_sc_hd__o211a_1 _26087_ (.A1(_02941_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08745_),
    .X(_08764_));
 sky130_fd_sc_hd__mux2_1 _26088_ (.A0(_08764_),
    .A1(net3028),
    .S(_08752_),
    .X(_08765_));
 sky130_fd_sc_hd__clkbuf_1 _26089_ (.A(_08765_),
    .X(_02697_));
 sky130_fd_sc_hd__o211a_1 _26090_ (.A1(_02946_),
    .A2(_08724_),
    .B1(_08725_),
    .C1(_08748_),
    .X(_08766_));
 sky130_fd_sc_hd__mux2_1 _26091_ (.A0(_08766_),
    .A1(net2515),
    .S(_08752_),
    .X(_08767_));
 sky130_fd_sc_hd__clkbuf_1 _26092_ (.A(_08767_),
    .X(_02698_));
 sky130_fd_sc_hd__buf_4 _26093_ (.A(_09125_),
    .X(_08768_));
 sky130_fd_sc_hd__o211a_1 _26094_ (.A1(_12169_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08727_),
    .X(_08769_));
 sky130_fd_sc_hd__mux2_1 _26095_ (.A0(_08769_),
    .A1(net2849),
    .S(_08752_),
    .X(_08770_));
 sky130_fd_sc_hd__clkbuf_1 _26096_ (.A(_08770_),
    .X(_02699_));
 sky130_fd_sc_hd__o211a_1 _26097_ (.A1(_12194_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08730_),
    .X(_08771_));
 sky130_fd_sc_hd__mux2_1 _26098_ (.A0(_08771_),
    .A1(net3484),
    .S(_08752_),
    .X(_08772_));
 sky130_fd_sc_hd__clkbuf_1 _26099_ (.A(_08772_),
    .X(_02700_));
 sky130_fd_sc_hd__o211a_1 _26100_ (.A1(_12202_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08733_),
    .X(_08773_));
 sky130_fd_sc_hd__mux2_1 _26101_ (.A0(_08773_),
    .A1(net2576),
    .S(_08752_),
    .X(_08774_));
 sky130_fd_sc_hd__clkbuf_1 _26102_ (.A(_08774_),
    .X(_02701_));
 sky130_fd_sc_hd__o211a_1 _26103_ (.A1(_12210_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08736_),
    .X(_08775_));
 sky130_fd_sc_hd__mux2_1 _26104_ (.A0(_08775_),
    .A1(net3201),
    .S(_08752_),
    .X(_08776_));
 sky130_fd_sc_hd__clkbuf_1 _26105_ (.A(_08776_),
    .X(_02702_));
 sky130_fd_sc_hd__o211a_1 _26106_ (.A1(_12218_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08739_),
    .X(_08777_));
 sky130_fd_sc_hd__mux2_1 _26107_ (.A0(_08777_),
    .A1(net2579),
    .S(_08752_),
    .X(_08778_));
 sky130_fd_sc_hd__clkbuf_1 _26108_ (.A(_08778_),
    .X(_02703_));
 sky130_fd_sc_hd__o211a_1 _26109_ (.A1(_12226_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08742_),
    .X(_08779_));
 sky130_fd_sc_hd__mux2_1 _26110_ (.A0(_08779_),
    .A1(net2865),
    .S(_08752_),
    .X(_08780_));
 sky130_fd_sc_hd__clkbuf_1 _26111_ (.A(_08780_),
    .X(_02704_));
 sky130_fd_sc_hd__o211a_1 _26112_ (.A1(_12234_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08745_),
    .X(_08781_));
 sky130_fd_sc_hd__mux2_1 _26113_ (.A0(_08781_),
    .A1(net3025),
    .S(_08752_),
    .X(_08782_));
 sky130_fd_sc_hd__clkbuf_1 _26114_ (.A(_08782_),
    .X(_02705_));
 sky130_fd_sc_hd__o211a_1 _26115_ (.A1(_12242_),
    .A2(_08726_),
    .B1(_08768_),
    .C1(_08748_),
    .X(_08783_));
 sky130_fd_sc_hd__mux2_1 _26116_ (.A0(_08783_),
    .A1(net2304),
    .S(_08752_),
    .X(_08784_));
 sky130_fd_sc_hd__clkbuf_1 _26117_ (.A(_08784_),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _26118_ (.A0(_07699_),
    .A1(net2879),
    .S(_12192_),
    .X(_08785_));
 sky130_fd_sc_hd__clkbuf_1 _26119_ (.A(_08785_),
    .X(_02707_));
 sky130_fd_sc_hd__mux2_1 _26120_ (.A0(_07703_),
    .A1(net2691),
    .S(_12192_),
    .X(_08786_));
 sky130_fd_sc_hd__clkbuf_1 _26121_ (.A(_08786_),
    .X(_02708_));
 sky130_fd_sc_hd__mux2_1 _26122_ (.A0(_07705_),
    .A1(net2294),
    .S(_12192_),
    .X(_08787_));
 sky130_fd_sc_hd__clkbuf_1 _26123_ (.A(_08787_),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_1 _26124_ (.A0(_07707_),
    .A1(net3416),
    .S(_12192_),
    .X(_08788_));
 sky130_fd_sc_hd__clkbuf_1 _26125_ (.A(_08788_),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _26126_ (.A0(_07709_),
    .A1(net3259),
    .S(_12192_),
    .X(_08789_));
 sky130_fd_sc_hd__clkbuf_1 _26127_ (.A(_08789_),
    .X(_02711_));
 sky130_fd_sc_hd__mux2_1 _26128_ (.A0(_07711_),
    .A1(net2904),
    .S(_12192_),
    .X(_08790_));
 sky130_fd_sc_hd__clkbuf_1 _26129_ (.A(_08790_),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _26130_ (.A0(_07713_),
    .A1(net3072),
    .S(_12192_),
    .X(_08791_));
 sky130_fd_sc_hd__clkbuf_1 _26131_ (.A(_08791_),
    .X(_02713_));
 sky130_fd_sc_hd__mux2_1 _26132_ (.A0(_07715_),
    .A1(net2670),
    .S(_12192_),
    .X(_08792_));
 sky130_fd_sc_hd__clkbuf_1 _26133_ (.A(_08792_),
    .X(_02714_));
 sky130_fd_sc_hd__o211a_1 _26134_ (.A1(_02850_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12186_),
    .X(_08793_));
 sky130_fd_sc_hd__clkbuf_8 _26135_ (.A(_12191_),
    .X(_08794_));
 sky130_fd_sc_hd__mux2_1 _26136_ (.A0(_08793_),
    .A1(net2802),
    .S(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__clkbuf_1 _26137_ (.A(_08795_),
    .X(_02715_));
 sky130_fd_sc_hd__o211a_1 _26138_ (.A1(_02860_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12199_),
    .X(_08796_));
 sky130_fd_sc_hd__mux2_1 _26139_ (.A0(_08796_),
    .A1(net3711),
    .S(_08794_),
    .X(_08797_));
 sky130_fd_sc_hd__clkbuf_1 _26140_ (.A(_08797_),
    .X(_02716_));
 sky130_fd_sc_hd__o211a_1 _26141_ (.A1(_02867_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12207_),
    .X(_08798_));
 sky130_fd_sc_hd__mux2_1 _26142_ (.A0(_08798_),
    .A1(net3168),
    .S(_08794_),
    .X(_08799_));
 sky130_fd_sc_hd__clkbuf_1 _26143_ (.A(_08799_),
    .X(_02717_));
 sky130_fd_sc_hd__o211a_1 _26144_ (.A1(_02874_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12215_),
    .X(_08800_));
 sky130_fd_sc_hd__mux2_1 _26145_ (.A0(_08800_),
    .A1(net2866),
    .S(_08794_),
    .X(_08801_));
 sky130_fd_sc_hd__clkbuf_1 _26146_ (.A(_08801_),
    .X(_02718_));
 sky130_fd_sc_hd__o211a_1 _26147_ (.A1(_02881_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12223_),
    .X(_08802_));
 sky130_fd_sc_hd__mux2_1 _26148_ (.A0(_08802_),
    .A1(net2311),
    .S(_08794_),
    .X(_08803_));
 sky130_fd_sc_hd__clkbuf_1 _26149_ (.A(_08803_),
    .X(_02719_));
 sky130_fd_sc_hd__o211a_1 _26150_ (.A1(_02888_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12231_),
    .X(_08804_));
 sky130_fd_sc_hd__mux2_1 _26151_ (.A0(_08804_),
    .A1(net2872),
    .S(_08794_),
    .X(_08805_));
 sky130_fd_sc_hd__clkbuf_1 _26152_ (.A(_08805_),
    .X(_02720_));
 sky130_fd_sc_hd__o211a_1 _26153_ (.A1(_02895_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12239_),
    .X(_08806_));
 sky130_fd_sc_hd__mux2_1 _26154_ (.A0(_08806_),
    .A1(net2871),
    .S(_08794_),
    .X(_08807_));
 sky130_fd_sc_hd__clkbuf_1 _26155_ (.A(_08807_),
    .X(_02721_));
 sky130_fd_sc_hd__o211a_1 _26156_ (.A1(_02902_),
    .A2(_12179_),
    .B1(_08768_),
    .C1(_12247_),
    .X(_08808_));
 sky130_fd_sc_hd__mux2_1 _26157_ (.A0(_08808_),
    .A1(net3614),
    .S(_08794_),
    .X(_08809_));
 sky130_fd_sc_hd__clkbuf_1 _26158_ (.A(_08809_),
    .X(_02722_));
 sky130_fd_sc_hd__o211a_1 _26159_ (.A1(_02910_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12186_),
    .X(_08810_));
 sky130_fd_sc_hd__mux2_1 _26160_ (.A0(_08810_),
    .A1(net3667),
    .S(_08794_),
    .X(_08811_));
 sky130_fd_sc_hd__clkbuf_1 _26161_ (.A(_08811_),
    .X(_02723_));
 sky130_fd_sc_hd__o211a_1 _26162_ (.A1(_02915_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12199_),
    .X(_08812_));
 sky130_fd_sc_hd__mux2_1 _26163_ (.A0(_08812_),
    .A1(net3600),
    .S(_08794_),
    .X(_08813_));
 sky130_fd_sc_hd__clkbuf_1 _26164_ (.A(_08813_),
    .X(_02724_));
 sky130_fd_sc_hd__o211a_1 _26165_ (.A1(_02920_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12207_),
    .X(_08814_));
 sky130_fd_sc_hd__mux2_1 _26166_ (.A0(_08814_),
    .A1(net3457),
    .S(_08794_),
    .X(_08815_));
 sky130_fd_sc_hd__clkbuf_1 _26167_ (.A(_08815_),
    .X(_02725_));
 sky130_fd_sc_hd__o211a_1 _26168_ (.A1(_02926_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12215_),
    .X(_08816_));
 sky130_fd_sc_hd__mux2_1 _26169_ (.A0(_08816_),
    .A1(net3127),
    .S(_08794_),
    .X(_08817_));
 sky130_fd_sc_hd__clkbuf_1 _26170_ (.A(_08817_),
    .X(_02726_));
 sky130_fd_sc_hd__o211a_1 _26171_ (.A1(_02931_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12223_),
    .X(_08818_));
 sky130_fd_sc_hd__mux2_1 _26172_ (.A0(_08818_),
    .A1(net3540),
    .S(_08794_),
    .X(_08819_));
 sky130_fd_sc_hd__clkbuf_1 _26173_ (.A(_08819_),
    .X(_02727_));
 sky130_fd_sc_hd__o211a_1 _26174_ (.A1(_02936_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12231_),
    .X(_08820_));
 sky130_fd_sc_hd__mux2_1 _26175_ (.A0(_08820_),
    .A1(net3531),
    .S(_08794_),
    .X(_08821_));
 sky130_fd_sc_hd__clkbuf_1 _26176_ (.A(_08821_),
    .X(_02728_));
 sky130_fd_sc_hd__o211a_1 _26177_ (.A1(_02941_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12239_),
    .X(_08822_));
 sky130_fd_sc_hd__mux2_1 _26178_ (.A0(_08822_),
    .A1(net3506),
    .S(_08794_),
    .X(_08823_));
 sky130_fd_sc_hd__clkbuf_1 _26179_ (.A(_08823_),
    .X(_02729_));
 sky130_fd_sc_hd__o211a_1 _26180_ (.A1(_02946_),
    .A2(_12182_),
    .B1(_12840_),
    .C1(_12247_),
    .X(_08824_));
 sky130_fd_sc_hd__mux2_1 _26181_ (.A0(_08824_),
    .A1(net3426),
    .S(_08794_),
    .X(_08825_));
 sky130_fd_sc_hd__clkbuf_1 _26182_ (.A(_08825_),
    .X(_02730_));
 sky130_fd_sc_hd__or2b_1 _26183_ (.A(net3885),
    .B_N(_09128_),
    .X(_08826_));
 sky130_fd_sc_hd__clkbuf_1 _26184_ (.A(net3886),
    .X(_02731_));
 sky130_fd_sc_hd__o21ai_1 _26185_ (.A1(_12188_),
    .A2(_09105_),
    .B1(_12328_),
    .Y(_08827_));
 sky130_fd_sc_hd__mux2_1 _26186_ (.A0(_09107_),
    .A1(net3998),
    .S(_08827_),
    .X(_08828_));
 sky130_fd_sc_hd__clkbuf_1 _26187_ (.A(net3999),
    .X(_02732_));
 sky130_fd_sc_hd__dfstp_1 _26188_ (.CLK(clknet_leaf_366_clk_i),
    .D(net1996),
    .SET_B(net141),
    .Q(\fb_read_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26189_ (.CLK(clknet_leaf_365_clk_i),
    .D(net3978),
    .RESET_B(net141),
    .Q(\fb_read_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26190_ (.CLK(clknet_leaf_366_clk_i),
    .D(net3973),
    .RESET_B(net141),
    .Q(\fb_read_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26191_ (.CLK(clknet_leaf_319_clk_i),
    .D(_00012_),
    .RESET_B(net259),
    .Q(\line_cache[319][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26192_ (.CLK(clknet_leaf_318_clk_i),
    .D(_00013_),
    .RESET_B(net259),
    .Q(\line_cache[319][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26193_ (.CLK(clknet_leaf_319_clk_i),
    .D(_00014_),
    .RESET_B(net259),
    .Q(\line_cache[319][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26194_ (.CLK(clknet_leaf_319_clk_i),
    .D(_00015_),
    .RESET_B(net259),
    .Q(\line_cache[319][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26195_ (.CLK(clknet_leaf_318_clk_i),
    .D(_00016_),
    .RESET_B(net263),
    .Q(\line_cache[319][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26196_ (.CLK(clknet_leaf_319_clk_i),
    .D(_00017_),
    .RESET_B(net259),
    .Q(\line_cache[319][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26197_ (.CLK(clknet_leaf_319_clk_i),
    .D(_00018_),
    .RESET_B(net263),
    .Q(\line_cache[319][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26198_ (.CLK(clknet_leaf_319_clk_i),
    .D(_00019_),
    .RESET_B(net263),
    .Q(\line_cache[319][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26199_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00020_),
    .RESET_B(net142),
    .Q(\res_v_active[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26200_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00021_),
    .RESET_B(net142),
    .Q(\res_v_active[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26201_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00022_),
    .RESET_B(net142),
    .Q(\res_v_active[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26202_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00023_),
    .RESET_B(net142),
    .Q(\res_v_active[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26203_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00024_),
    .RESET_B(net142),
    .Q(\res_v_active[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26204_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00025_),
    .RESET_B(net142),
    .Q(\res_v_active[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26205_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00026_),
    .RESET_B(net142),
    .Q(\res_v_active[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26206_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00027_),
    .RESET_B(net142),
    .Q(\res_v_active[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26207_ (.CLK(clknet_leaf_339_clk_i),
    .D(_00028_),
    .RESET_B(net171),
    .Q(\line_cache_idx[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26208_ (.CLK(clknet_leaf_339_clk_i),
    .D(net3922),
    .RESET_B(net171),
    .Q(\line_cache_idx[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26209_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00030_),
    .RESET_B(net176),
    .Q(\line_cache_idx[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26210_ (.CLK(clknet_leaf_33_clk_i),
    .D(net3382),
    .RESET_B(net179),
    .Q(\line_cache_idx[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26211_ (.CLK(clknet_leaf_328_clk_i),
    .D(_00032_),
    .RESET_B(net183),
    .Q(\line_cache_idx[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26212_ (.CLK(clknet_leaf_39_clk_i),
    .D(net3914),
    .RESET_B(net183),
    .Q(\line_cache_idx[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26213_ (.CLK(clknet_leaf_328_clk_i),
    .D(_00034_),
    .RESET_B(net181),
    .Q(\line_cache_idx[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26214_ (.CLK(clknet_leaf_328_clk_i),
    .D(_00035_),
    .RESET_B(net181),
    .Q(\line_cache_idx[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26215_ (.CLK(clknet_leaf_296_clk_i),
    .D(net2562),
    .RESET_B(net251),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _26216_ (.CLK(clknet_leaf_296_clk_i),
    .D(net3901),
    .RESET_B(net251),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _26217_ (.CLK(clknet_leaf_295_clk_i),
    .D(net3558),
    .RESET_B(net251),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _26218_ (.CLK(clknet_leaf_295_clk_i),
    .D(net3765),
    .RESET_B(net253),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _26219_ (.CLK(clknet_leaf_295_clk_i),
    .D(net3856),
    .RESET_B(net251),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _26220_ (.CLK(clknet_leaf_294_clk_i),
    .D(_00041_),
    .RESET_B(net253),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _26221_ (.CLK(clknet_leaf_294_clk_i),
    .D(net3625),
    .RESET_B(net253),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _26222_ (.CLK(clknet_leaf_294_clk_i),
    .D(net2751),
    .RESET_B(net253),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _26223_ (.CLK(clknet_leaf_294_clk_i),
    .D(net3619),
    .RESET_B(net253),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _26224_ (.CLK(clknet_leaf_293_clk_i),
    .D(net3769),
    .RESET_B(net253),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _26225_ (.CLK(clknet_leaf_294_clk_i),
    .D(net3822),
    .RESET_B(net269),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _26226_ (.CLK(clknet_leaf_281_clk_i),
    .D(net3498),
    .RESET_B(net269),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _26227_ (.CLK(clknet_leaf_281_clk_i),
    .D(net3791),
    .RESET_B(net269),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_2 _26228_ (.CLK(clknet_leaf_281_clk_i),
    .D(net3495),
    .RESET_B(net269),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _26229_ (.CLK(clknet_leaf_280_clk_i),
    .D(net3793),
    .RESET_B(net269),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _26230_ (.CLK(clknet_leaf_280_clk_i),
    .D(net3661),
    .RESET_B(net269),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _26231_ (.CLK(clknet_leaf_280_clk_i),
    .D(net3848),
    .RESET_B(net271),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _26232_ (.CLK(clknet_leaf_280_clk_i),
    .D(net2010),
    .RESET_B(net271),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _26233_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00054_),
    .RESET_B(net271),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 _26234_ (.CLK(clknet_leaf_279_clk_i),
    .D(net3017),
    .RESET_B(net271),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_2 _26235_ (.CLK(clknet_leaf_279_clk_i),
    .D(net3843),
    .RESET_B(net271),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _26236_ (.CLK(clknet_leaf_279_clk_i),
    .D(net2022),
    .RESET_B(net271),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _26237_ (.CLK(clknet_leaf_279_clk_i),
    .D(net3862),
    .RESET_B(net277),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _26238_ (.CLK(clknet_leaf_279_clk_i),
    .D(net3608),
    .RESET_B(net277),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _26239_ (.CLK(clknet_leaf_276_clk_i),
    .D(net3951),
    .RESET_B(net277),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _26240_ (.CLK(clknet_leaf_276_clk_i),
    .D(net2018),
    .RESET_B(net277),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_1 _26241_ (.CLK(clknet_leaf_275_clk_i),
    .D(_00062_),
    .RESET_B(net277),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_1 _26242_ (.CLK(clknet_leaf_276_clk_i),
    .D(net2008),
    .RESET_B(net277),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _26243_ (.CLK(clknet_leaf_275_clk_i),
    .D(net3957),
    .RESET_B(net277),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_1 _26244_ (.CLK(clknet_leaf_275_clk_i),
    .D(net3963),
    .RESET_B(net277),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _26245_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00066_),
    .RESET_B(net137),
    .Q(\prescaler[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26246_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00067_),
    .RESET_B(net137),
    .Q(\prescaler[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26247_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00068_),
    .RESET_B(net137),
    .Q(\prescaler[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26248_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00069_),
    .RESET_B(net137),
    .Q(\prescaler[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26249_ (.CLK(clknet_leaf_367_clk_i),
    .D(_00070_),
    .RESET_B(net140),
    .Q(\resolution[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26250_ (.CLK(clknet_leaf_367_clk_i),
    .D(_00071_),
    .RESET_B(net140),
    .Q(\resolution[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26251_ (.CLK(clknet_leaf_367_clk_i),
    .D(_00072_),
    .RESET_B(net140),
    .Q(\resolution[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26252_ (.CLK(clknet_leaf_367_clk_i),
    .D(_00073_),
    .RESET_B(net140),
    .Q(\resolution[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26253_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00074_),
    .RESET_B(net138),
    .Q(\base_h_active[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26254_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00075_),
    .RESET_B(net138),
    .Q(\base_h_active[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26255_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00076_),
    .RESET_B(net138),
    .Q(\base_h_active[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26256_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00077_),
    .RESET_B(net139),
    .Q(\base_h_active[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26257_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00078_),
    .RESET_B(net137),
    .Q(\base_h_active[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26258_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00079_),
    .RESET_B(net137),
    .Q(\base_h_active[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26259_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00080_),
    .RESET_B(net139),
    .Q(\base_h_active[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26260_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00081_),
    .RESET_B(net139),
    .Q(\base_h_active[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26261_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00082_),
    .RESET_B(net139),
    .Q(\base_h_active[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26262_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00083_),
    .RESET_B(net139),
    .Q(\base_h_active[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26263_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00084_),
    .RESET_B(net138),
    .Q(\base_h_fporch[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26264_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00085_),
    .RESET_B(net138),
    .Q(\base_h_fporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26265_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00086_),
    .RESET_B(net138),
    .Q(\base_h_fporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26266_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00087_),
    .RESET_B(net138),
    .Q(\base_h_fporch[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26267_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00088_),
    .RESET_B(net137),
    .Q(\base_h_fporch[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26268_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00089_),
    .RESET_B(net138),
    .Q(\base_h_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26269_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00090_),
    .RESET_B(net138),
    .Q(\base_h_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26270_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00091_),
    .RESET_B(net138),
    .Q(\base_h_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26271_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00092_),
    .RESET_B(net138),
    .Q(\base_h_sync[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26272_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00093_),
    .RESET_B(net137),
    .Q(\base_h_sync[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26273_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00094_),
    .RESET_B(net137),
    .Q(\base_h_sync[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26274_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00095_),
    .RESET_B(net137),
    .Q(\base_h_sync[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26275_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00096_),
    .RESET_B(net138),
    .Q(\base_h_bporch[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26276_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00097_),
    .RESET_B(net138),
    .Q(\base_h_bporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26277_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00098_),
    .RESET_B(net138),
    .Q(\base_h_bporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26278_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00099_),
    .RESET_B(net138),
    .Q(\base_h_bporch[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26279_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00100_),
    .RESET_B(net137),
    .Q(\base_h_bporch[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26280_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00101_),
    .RESET_B(net137),
    .Q(\base_h_bporch[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26281_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00102_),
    .RESET_B(net137),
    .Q(\base_h_bporch[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26282_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00103_),
    .RESET_B(net150),
    .Q(\base_v_active[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26283_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00104_),
    .RESET_B(net150),
    .Q(\base_v_active[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26284_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00105_),
    .RESET_B(net150),
    .Q(\base_v_active[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26285_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00106_),
    .RESET_B(net150),
    .Q(\base_v_active[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26286_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00107_),
    .RESET_B(net150),
    .Q(\base_v_active[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26287_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00108_),
    .RESET_B(net150),
    .Q(\base_v_active[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26288_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00109_),
    .RESET_B(net150),
    .Q(\base_v_active[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26289_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00110_),
    .RESET_B(net150),
    .Q(\base_v_active[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26290_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00111_),
    .RESET_B(net138),
    .Q(\base_v_active[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26291_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00112_),
    .RESET_B(net150),
    .Q(\base_v_fporch[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26292_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00113_),
    .RESET_B(net147),
    .Q(\base_v_fporch[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26293_ (.CLK(clknet_5_2__leaf_clk_i),
    .D(_00114_),
    .RESET_B(net150),
    .Q(\base_v_fporch[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26294_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00115_),
    .RESET_B(net147),
    .Q(\base_v_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26295_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00116_),
    .RESET_B(net147),
    .Q(\base_v_sync[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26296_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00117_),
    .RESET_B(net147),
    .Q(\base_v_sync[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26297_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00118_),
    .RESET_B(net147),
    .Q(\base_v_bporch[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26298_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00119_),
    .RESET_B(net147),
    .Q(\base_v_bporch[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26299_ (.CLK(clknet_leaf_67_clk_i),
    .D(_00120_),
    .RESET_B(net186),
    .Q(\base_v_bporch[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26300_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00121_),
    .RESET_B(net147),
    .Q(\base_v_bporch[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26301_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00000_),
    .RESET_B(net137),
    .Q(\prescaler_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26302_ (.CLK(clknet_leaf_371_clk_i),
    .D(_00001_),
    .RESET_B(net137),
    .Q(\prescaler_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26303_ (.CLK(clknet_leaf_370_clk_i),
    .D(_00002_),
    .RESET_B(net137),
    .Q(\prescaler_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26304_ (.CLK(clknet_leaf_370_clk_i),
    .D(_00003_),
    .RESET_B(net146),
    .Q(\prescaler_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26305_ (.CLK(clknet_leaf_370_clk_i),
    .D(_00004_),
    .RESET_B(net146),
    .Q(\prescaler_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26306_ (.CLK(clknet_leaf_370_clk_i),
    .D(_00005_),
    .RESET_B(net146),
    .Q(\prescaler_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26307_ (.CLK(clknet_leaf_370_clk_i),
    .D(_00006_),
    .RESET_B(net146),
    .Q(\prescaler_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26308_ (.CLK(clknet_leaf_367_clk_i),
    .D(_00007_),
    .RESET_B(net140),
    .Q(\prescaler_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26309_ (.CLK(clknet_leaf_367_clk_i),
    .D(_00008_),
    .RESET_B(net140),
    .Q(\prescaler_counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26310_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00122_),
    .RESET_B(net142),
    .Q(\res_h_active[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26311_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00123_),
    .RESET_B(net142),
    .Q(\res_h_active[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26312_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00124_),
    .RESET_B(net151),
    .Q(\res_h_active[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26313_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00125_),
    .RESET_B(net151),
    .Q(\res_h_active[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26314_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00126_),
    .RESET_B(net151),
    .Q(\res_h_active[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26315_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00127_),
    .RESET_B(net151),
    .Q(\res_h_active[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26316_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00128_),
    .RESET_B(net151),
    .Q(\res_h_active[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26317_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00129_),
    .RESET_B(net151),
    .Q(\res_h_active[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26318_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00130_),
    .RESET_B(net151),
    .Q(\res_h_active[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26319_ (.CLK(clknet_leaf_5_clk_i),
    .D(net1986),
    .RESET_B(net142),
    .Q(\base_h_counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26320_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00132_),
    .RESET_B(net139),
    .Q(\base_h_counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26321_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00133_),
    .RESET_B(net139),
    .Q(\base_h_counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26322_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00134_),
    .RESET_B(net139),
    .Q(\base_h_counter[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26323_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00135_),
    .RESET_B(net139),
    .Q(\base_h_counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26324_ (.CLK(clknet_leaf_1_clk_i),
    .D(net3993),
    .RESET_B(net139),
    .Q(\base_h_counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26325_ (.CLK(clknet_5_1__leaf_clk_i),
    .D(_00137_),
    .RESET_B(net140),
    .Q(\base_h_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26326_ (.CLK(clknet_leaf_368_clk_i),
    .D(net3969),
    .RESET_B(net140),
    .Q(\base_h_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26327_ (.CLK(clknet_leaf_368_clk_i),
    .D(net3960),
    .RESET_B(net140),
    .Q(\base_h_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26328_ (.CLK(clknet_leaf_368_clk_i),
    .D(net3948),
    .RESET_B(net140),
    .Q(\base_h_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26329_ (.CLK(clknet_leaf_11_clk_i),
    .D(net2027),
    .RESET_B(net151),
    .Q(\base_v_counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26330_ (.CLK(clknet_leaf_11_clk_i),
    .D(net3802),
    .RESET_B(net150),
    .Q(\base_v_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26331_ (.CLK(clknet_leaf_11_clk_i),
    .D(net2013),
    .RESET_B(net151),
    .Q(\base_v_counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26332_ (.CLK(clknet_leaf_11_clk_i),
    .D(net3786),
    .RESET_B(net151),
    .Q(\base_v_counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26333_ (.CLK(clknet_leaf_10_clk_i),
    .D(net3799),
    .RESET_B(net151),
    .Q(\base_v_counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26334_ (.CLK(clknet_leaf_10_clk_i),
    .D(net3819),
    .RESET_B(net151),
    .Q(\base_v_counter[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26335_ (.CLK(clknet_leaf_10_clk_i),
    .D(net3814),
    .RESET_B(net151),
    .Q(\base_v_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26336_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00148_),
    .RESET_B(net142),
    .Q(\base_v_counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26337_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00149_),
    .RESET_B(net142),
    .Q(\base_v_counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26338_ (.CLK(clknet_leaf_4_clk_i),
    .D(net3715),
    .RESET_B(net139),
    .Q(\base_v_counter[9] ));
 sky130_fd_sc_hd__dfrtp_4 _26339_ (.CLK(clknet_leaf_339_clk_i),
    .D(net3774),
    .RESET_B(net171),
    .Q(\res_h_counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26340_ (.CLK(clknet_leaf_331_clk_i),
    .D(net3868),
    .RESET_B(net181),
    .Q(\res_h_counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26341_ (.CLK(clknet_leaf_332_clk_i),
    .D(net3746),
    .RESET_B(net181),
    .Q(\res_h_counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26342_ (.CLK(clknet_leaf_331_clk_i),
    .D(net3639),
    .RESET_B(net181),
    .Q(\res_h_counter[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26343_ (.CLK(clknet_leaf_332_clk_i),
    .D(net3944),
    .RESET_B(net181),
    .Q(\res_h_counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26344_ (.CLK(clknet_leaf_332_clk_i),
    .D(net3903),
    .RESET_B(net181),
    .Q(\res_h_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26345_ (.CLK(clknet_leaf_332_clk_i),
    .D(net1998),
    .RESET_B(net181),
    .Q(\res_h_counter[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26346_ (.CLK(clknet_leaf_329_clk_i),
    .D(net3916),
    .RESET_B(net181),
    .Q(\res_h_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26347_ (.CLK(clknet_leaf_332_clk_i),
    .D(_00159_),
    .RESET_B(net181),
    .Q(\res_h_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26348_ (.CLK(clknet_leaf_339_clk_i),
    .D(net1960),
    .RESET_B(net171),
    .Q(\res_h_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26349_ (.CLK(clknet_leaf_364_clk_i),
    .D(net3830),
    .RESET_B(net140),
    .Q(\res_v_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26350_ (.CLK(clknet_leaf_364_clk_i),
    .D(net2004),
    .RESET_B(net142),
    .Q(\res_v_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26351_ (.CLK(clknet_leaf_5_clk_i),
    .D(net3805),
    .RESET_B(net142),
    .Q(\res_v_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26352_ (.CLK(clknet_leaf_363_clk_i),
    .D(net3750),
    .RESET_B(net142),
    .Q(\res_v_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26353_ (.CLK(clknet_leaf_364_clk_i),
    .D(net2498),
    .RESET_B(net140),
    .Q(\res_v_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26354_ (.CLK(clknet_leaf_364_clk_i),
    .D(net3778),
    .RESET_B(net143),
    .Q(\res_v_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26355_ (.CLK(clknet_leaf_364_clk_i),
    .D(net3452),
    .RESET_B(net141),
    .Q(\res_v_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26356_ (.CLK(clknet_leaf_364_clk_i),
    .D(net3837),
    .RESET_B(net141),
    .Q(\res_v_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26357_ (.CLK(clknet_leaf_364_clk_i),
    .D(net2029),
    .RESET_B(net140),
    .Q(\res_v_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26358_ (.CLK(clknet_leaf_364_clk_i),
    .D(net2058),
    .RESET_B(net140),
    .Q(\res_v_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26359_ (.CLK(clknet_leaf_366_clk_i),
    .D(net2016),
    .RESET_B(net141),
    .Q(\pixel_double_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26360_ (.CLK(clknet_leaf_367_clk_i),
    .D(net2001),
    .RESET_B(net140),
    .Q(\pixel_double_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26361_ (.CLK(clknet_leaf_367_clk_i),
    .D(net1942),
    .RESET_B(net140),
    .Q(\pixel_double_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26362_ (.CLK(clknet_leaf_368_clk_i),
    .D(net1864),
    .RESET_B(net145),
    .Q(\pixel_double_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26363_ (.CLK(clknet_leaf_366_clk_i),
    .D(net2112),
    .RESET_B(net141),
    .Q(\line_double_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26364_ (.CLK(clknet_leaf_366_clk_i),
    .D(net2798),
    .RESET_B(net141),
    .Q(\line_double_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26365_ (.CLK(clknet_leaf_366_clk_i),
    .D(net1993),
    .RESET_B(net141),
    .Q(\line_double_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26366_ (.CLK(clknet_leaf_367_clk_i),
    .D(net2006),
    .RESET_B(net141),
    .Q(\line_double_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26367_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00179_),
    .RESET_B(net263),
    .Q(\line_cache[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26368_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00180_),
    .RESET_B(net263),
    .Q(\line_cache[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26369_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00181_),
    .RESET_B(net265),
    .Q(\line_cache[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26370_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00182_),
    .RESET_B(net263),
    .Q(\line_cache[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26371_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00183_),
    .RESET_B(net265),
    .Q(\line_cache[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26372_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00184_),
    .RESET_B(net307),
    .Q(\line_cache[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26373_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00185_),
    .RESET_B(net307),
    .Q(\line_cache[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26374_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00186_),
    .RESET_B(net307),
    .Q(\line_cache[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26375_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00187_),
    .RESET_B(net265),
    .Q(\line_cache[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26376_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00188_),
    .RESET_B(net265),
    .Q(\line_cache[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26377_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00189_),
    .RESET_B(net265),
    .Q(\line_cache[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26378_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00190_),
    .RESET_B(net266),
    .Q(\line_cache[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26379_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00191_),
    .RESET_B(net266),
    .Q(\line_cache[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26380_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00192_),
    .RESET_B(net267),
    .Q(\line_cache[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26381_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00193_),
    .RESET_B(net309),
    .Q(\line_cache[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26382_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00194_),
    .RESET_B(net309),
    .Q(\line_cache[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26383_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00195_),
    .RESET_B(net267),
    .Q(\line_cache[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26384_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00196_),
    .RESET_B(net267),
    .Q(\line_cache[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26385_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00197_),
    .RESET_B(net307),
    .Q(\line_cache[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26386_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00198_),
    .RESET_B(net267),
    .Q(\line_cache[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26387_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00199_),
    .RESET_B(net267),
    .Q(\line_cache[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26388_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00200_),
    .RESET_B(net267),
    .Q(\line_cache[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26389_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00201_),
    .RESET_B(net309),
    .Q(\line_cache[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26390_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00202_),
    .RESET_B(net309),
    .Q(\line_cache[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26391_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00203_),
    .RESET_B(net265),
    .Q(\line_cache[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26392_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00204_),
    .RESET_B(net265),
    .Q(\line_cache[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26393_ (.CLK(clknet_leaf_231_clk_i),
    .D(_00205_),
    .RESET_B(net267),
    .Q(\line_cache[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26394_ (.CLK(clknet_leaf_232_clk_i),
    .D(_00206_),
    .RESET_B(net267),
    .Q(\line_cache[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26395_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00207_),
    .RESET_B(net266),
    .Q(\line_cache[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26396_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00208_),
    .RESET_B(net266),
    .Q(\line_cache[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26397_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00209_),
    .RESET_B(net266),
    .Q(\line_cache[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26398_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00210_),
    .RESET_B(net266),
    .Q(\line_cache[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26399_ (.CLK(clknet_leaf_230_clk_i),
    .D(_00211_),
    .RESET_B(net265),
    .Q(\line_cache[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26400_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00212_),
    .RESET_B(net265),
    .Q(\line_cache[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26401_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00213_),
    .RESET_B(net265),
    .Q(\line_cache[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26402_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00214_),
    .RESET_B(net266),
    .Q(\line_cache[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26403_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00215_),
    .RESET_B(net266),
    .Q(\line_cache[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26404_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00216_),
    .RESET_B(net266),
    .Q(\line_cache[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26405_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00217_),
    .RESET_B(net266),
    .Q(\line_cache[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26406_ (.CLK(clknet_leaf_235_clk_i),
    .D(_00218_),
    .RESET_B(net266),
    .Q(\line_cache[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26407_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00219_),
    .RESET_B(net266),
    .Q(\line_cache[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26408_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00220_),
    .RESET_B(net266),
    .Q(\line_cache[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26409_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00221_),
    .RESET_B(net288),
    .Q(\line_cache[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26410_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00222_),
    .RESET_B(net288),
    .Q(\line_cache[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26411_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00223_),
    .RESET_B(net288),
    .Q(\line_cache[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26412_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00224_),
    .RESET_B(net288),
    .Q(\line_cache[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26413_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00225_),
    .RESET_B(net288),
    .Q(\line_cache[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26414_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00226_),
    .RESET_B(net288),
    .Q(\line_cache[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26415_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00227_),
    .RESET_B(net266),
    .Q(\line_cache[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26416_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00228_),
    .RESET_B(net266),
    .Q(\line_cache[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26417_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00229_),
    .RESET_B(net288),
    .Q(\line_cache[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26418_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00230_),
    .RESET_B(net288),
    .Q(\line_cache[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26419_ (.CLK(clknet_leaf_234_clk_i),
    .D(_00231_),
    .RESET_B(net266),
    .Q(\line_cache[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26420_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00232_),
    .RESET_B(net288),
    .Q(\line_cache[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26421_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00233_),
    .RESET_B(net288),
    .Q(\line_cache[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26422_ (.CLK(clknet_leaf_245_clk_i),
    .D(_00234_),
    .RESET_B(net289),
    .Q(\line_cache[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26423_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00235_),
    .RESET_B(net288),
    .Q(\line_cache[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26424_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00236_),
    .RESET_B(net288),
    .Q(\line_cache[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26425_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00237_),
    .RESET_B(net288),
    .Q(\line_cache[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26426_ (.CLK(clknet_leaf_244_clk_i),
    .D(_00238_),
    .RESET_B(net288),
    .Q(\line_cache[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26427_ (.CLK(clknet_leaf_245_clk_i),
    .D(_00239_),
    .RESET_B(net289),
    .Q(\line_cache[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26428_ (.CLK(clknet_leaf_245_clk_i),
    .D(_00240_),
    .RESET_B(net288),
    .Q(\line_cache[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26429_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00241_),
    .RESET_B(net290),
    .Q(\line_cache[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26430_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00242_),
    .RESET_B(net288),
    .Q(\line_cache[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26431_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00243_),
    .RESET_B(net290),
    .Q(\line_cache[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26432_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00244_),
    .RESET_B(net290),
    .Q(\line_cache[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26433_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00245_),
    .RESET_B(net290),
    .Q(\line_cache[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26434_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00246_),
    .RESET_B(net290),
    .Q(\line_cache[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26435_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00247_),
    .RESET_B(net290),
    .Q(\line_cache[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26436_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00248_),
    .RESET_B(net290),
    .Q(\line_cache[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26437_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00249_),
    .RESET_B(net290),
    .Q(\line_cache[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26438_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00250_),
    .RESET_B(net290),
    .Q(\line_cache[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26439_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00251_),
    .RESET_B(net296),
    .Q(\line_cache[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26440_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00252_),
    .RESET_B(net296),
    .Q(\line_cache[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26441_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00253_),
    .RESET_B(net297),
    .Q(\line_cache[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26442_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00254_),
    .RESET_B(net296),
    .Q(\line_cache[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26443_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00255_),
    .RESET_B(net297),
    .Q(\line_cache[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26444_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00256_),
    .RESET_B(net296),
    .Q(\line_cache[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26445_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00257_),
    .RESET_B(net297),
    .Q(\line_cache[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26446_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00258_),
    .RESET_B(net298),
    .Q(\line_cache[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26447_ (.CLK(clknet_leaf_249_clk_i),
    .D(_00259_),
    .RESET_B(net290),
    .Q(\line_cache[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26448_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00260_),
    .RESET_B(net296),
    .Q(\line_cache[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26449_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00261_),
    .RESET_B(net297),
    .Q(\line_cache[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26450_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00262_),
    .RESET_B(net296),
    .Q(\line_cache[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26451_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00263_),
    .RESET_B(net298),
    .Q(\line_cache[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26452_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00264_),
    .RESET_B(net296),
    .Q(\line_cache[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26453_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00265_),
    .RESET_B(net298),
    .Q(\line_cache[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26454_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00266_),
    .RESET_B(net297),
    .Q(\line_cache[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26455_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00267_),
    .RESET_B(net296),
    .Q(\line_cache[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26456_ (.CLK(clknet_leaf_251_clk_i),
    .D(_00268_),
    .RESET_B(net296),
    .Q(\line_cache[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26457_ (.CLK(clknet_leaf_252_clk_i),
    .D(_00269_),
    .RESET_B(net298),
    .Q(\line_cache[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26458_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00270_),
    .RESET_B(net299),
    .Q(\line_cache[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26459_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00271_),
    .RESET_B(net298),
    .Q(\line_cache[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26460_ (.CLK(clknet_leaf_252_clk_i),
    .D(_00272_),
    .RESET_B(net299),
    .Q(\line_cache[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26461_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00273_),
    .RESET_B(net298),
    .Q(\line_cache[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26462_ (.CLK(clknet_leaf_252_clk_i),
    .D(_00274_),
    .RESET_B(net299),
    .Q(\line_cache[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26463_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00275_),
    .RESET_B(net335),
    .Q(\line_cache[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26464_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00276_),
    .RESET_B(net290),
    .Q(\line_cache[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26465_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00277_),
    .RESET_B(net290),
    .Q(\line_cache[12][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26466_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00278_),
    .RESET_B(net290),
    .Q(\line_cache[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26467_ (.CLK(clknet_leaf_252_clk_i),
    .D(_00279_),
    .RESET_B(net299),
    .Q(\line_cache[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26468_ (.CLK(clknet_leaf_252_clk_i),
    .D(_00280_),
    .RESET_B(net299),
    .Q(\line_cache[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26469_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00281_),
    .RESET_B(net298),
    .Q(\line_cache[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26470_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00282_),
    .RESET_B(net335),
    .Q(\line_cache[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26471_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00283_),
    .RESET_B(net291),
    .Q(\line_cache[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26472_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00284_),
    .RESET_B(net291),
    .Q(\line_cache[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26473_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00285_),
    .RESET_B(net289),
    .Q(\line_cache[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26474_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00286_),
    .RESET_B(net291),
    .Q(\line_cache[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26475_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00287_),
    .RESET_B(net329),
    .Q(\line_cache[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26476_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00288_),
    .RESET_B(net329),
    .Q(\line_cache[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26477_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00289_),
    .RESET_B(net328),
    .Q(\line_cache[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26478_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00290_),
    .RESET_B(net328),
    .Q(\line_cache[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26479_ (.CLK(clknet_leaf_248_clk_i),
    .D(_00291_),
    .RESET_B(net291),
    .Q(\line_cache[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26480_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00292_),
    .RESET_B(net291),
    .Q(\line_cache[14][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26481_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00293_),
    .RESET_B(net289),
    .Q(\line_cache[14][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26482_ (.CLK(clknet_leaf_247_clk_i),
    .D(_00294_),
    .RESET_B(net291),
    .Q(\line_cache[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26483_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00295_),
    .RESET_B(net329),
    .Q(\line_cache[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26484_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00296_),
    .RESET_B(net329),
    .Q(\line_cache[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26485_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00297_),
    .RESET_B(net328),
    .Q(\line_cache[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26486_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00298_),
    .RESET_B(net328),
    .Q(\line_cache[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26487_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00299_),
    .RESET_B(net267),
    .Q(\line_cache[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26488_ (.CLK(clknet_leaf_245_clk_i),
    .D(_00300_),
    .RESET_B(net289),
    .Q(\line_cache[15][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26489_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00301_),
    .RESET_B(net328),
    .Q(\line_cache[15][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26490_ (.CLK(clknet_leaf_246_clk_i),
    .D(_00302_),
    .RESET_B(net289),
    .Q(\line_cache[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26491_ (.CLK(clknet_leaf_233_clk_i),
    .D(_00303_),
    .RESET_B(net267),
    .Q(\line_cache[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26492_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00304_),
    .RESET_B(net309),
    .Q(\line_cache[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26493_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00305_),
    .RESET_B(net309),
    .Q(\line_cache[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26494_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00306_),
    .RESET_B(net328),
    .Q(\line_cache[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26495_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00307_),
    .RESET_B(net284),
    .Q(\line_cache[16][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26496_ (.CLK(clknet_leaf_265_clk_i),
    .D(_00308_),
    .RESET_B(net274),
    .Q(\line_cache[16][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26497_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00309_),
    .RESET_B(net284),
    .Q(\line_cache[16][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26498_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00310_),
    .RESET_B(net274),
    .Q(\line_cache[16][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26499_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00311_),
    .RESET_B(net274),
    .Q(\line_cache[16][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26500_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00312_),
    .RESET_B(net285),
    .Q(\line_cache[16][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26501_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00313_),
    .RESET_B(net285),
    .Q(\line_cache[16][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26502_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00314_),
    .RESET_B(net284),
    .Q(\line_cache[16][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26503_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00315_),
    .RESET_B(net273),
    .Q(\line_cache[17][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26504_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00316_),
    .RESET_B(net274),
    .Q(\line_cache[17][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26505_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00317_),
    .RESET_B(net284),
    .Q(\line_cache[17][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26506_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00318_),
    .RESET_B(net275),
    .Q(\line_cache[17][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26507_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00319_),
    .RESET_B(net275),
    .Q(\line_cache[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26508_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00320_),
    .RESET_B(net285),
    .Q(\line_cache[17][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26509_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00321_),
    .RESET_B(net285),
    .Q(\line_cache[17][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26510_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00322_),
    .RESET_B(net284),
    .Q(\line_cache[17][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26511_ (.CLK(clknet_leaf_286_clk_i),
    .D(_00323_),
    .RESET_B(net273),
    .Q(\line_cache[18][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26512_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00324_),
    .RESET_B(net273),
    .Q(\line_cache[18][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26513_ (.CLK(clknet_leaf_287_clk_i),
    .D(_00325_),
    .RESET_B(net273),
    .Q(\line_cache[18][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26514_ (.CLK(clknet_leaf_266_clk_i),
    .D(_00326_),
    .RESET_B(net275),
    .Q(\line_cache[18][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26515_ (.CLK(clknet_leaf_266_clk_i),
    .D(_00327_),
    .RESET_B(net274),
    .Q(\line_cache[18][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26516_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00328_),
    .RESET_B(net285),
    .Q(\line_cache[18][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26517_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00329_),
    .RESET_B(net275),
    .Q(\line_cache[18][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26518_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00330_),
    .RESET_B(net273),
    .Q(\line_cache[18][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26519_ (.CLK(clknet_leaf_286_clk_i),
    .D(_00331_),
    .RESET_B(net276),
    .Q(\line_cache[19][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26520_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00332_),
    .RESET_B(net276),
    .Q(\line_cache[19][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26521_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00333_),
    .RESET_B(net284),
    .Q(\line_cache[19][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26522_ (.CLK(clknet_leaf_284_clk_i),
    .D(_00334_),
    .RESET_B(net274),
    .Q(\line_cache[19][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26523_ (.CLK(clknet_leaf_265_clk_i),
    .D(_00335_),
    .RESET_B(net275),
    .Q(\line_cache[19][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26524_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00336_),
    .RESET_B(net285),
    .Q(\line_cache[19][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26525_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00337_),
    .RESET_B(net285),
    .Q(\line_cache[19][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26526_ (.CLK(clknet_leaf_264_clk_i),
    .D(_00338_),
    .RESET_B(net276),
    .Q(\line_cache[19][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26527_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00339_),
    .RESET_B(net284),
    .Q(\line_cache[20][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26528_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00340_),
    .RESET_B(net285),
    .Q(\line_cache[20][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26529_ (.CLK(clknet_leaf_237_clk_i),
    .D(_00341_),
    .RESET_B(net264),
    .Q(\line_cache[20][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26530_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00342_),
    .RESET_B(net285),
    .Q(\line_cache[20][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26531_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00343_),
    .RESET_B(net286),
    .Q(\line_cache[20][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26532_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00344_),
    .RESET_B(net286),
    .Q(\line_cache[20][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26533_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00345_),
    .RESET_B(net284),
    .Q(\line_cache[20][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26534_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00346_),
    .RESET_B(net284),
    .Q(\line_cache[20][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26535_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00347_),
    .RESET_B(net284),
    .Q(\line_cache[21][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26536_ (.CLK(clknet_leaf_241_clk_i),
    .D(_00348_),
    .RESET_B(net286),
    .Q(\line_cache[21][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26537_ (.CLK(clknet_leaf_237_clk_i),
    .D(_00349_),
    .RESET_B(net264),
    .Q(\line_cache[21][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26538_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00350_),
    .RESET_B(net285),
    .Q(\line_cache[21][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26539_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00351_),
    .RESET_B(net286),
    .Q(\line_cache[21][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26540_ (.CLK(clknet_leaf_241_clk_i),
    .D(_00352_),
    .RESET_B(net286),
    .Q(\line_cache[21][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26541_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00353_),
    .RESET_B(net284),
    .Q(\line_cache[21][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26542_ (.CLK(clknet_leaf_237_clk_i),
    .D(_00354_),
    .RESET_B(net284),
    .Q(\line_cache[21][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26543_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00355_),
    .RESET_B(net287),
    .Q(\line_cache[22][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26544_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00356_),
    .RESET_B(net286),
    .Q(\line_cache[22][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26545_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00357_),
    .RESET_B(net264),
    .Q(\line_cache[22][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26546_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00358_),
    .RESET_B(net290),
    .Q(\line_cache[22][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26547_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00359_),
    .RESET_B(net290),
    .Q(\line_cache[22][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26548_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00360_),
    .RESET_B(net287),
    .Q(\line_cache[22][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26549_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00361_),
    .RESET_B(net287),
    .Q(\line_cache[22][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26550_ (.CLK(clknet_leaf_237_clk_i),
    .D(_00362_),
    .RESET_B(net287),
    .Q(\line_cache[22][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26551_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00363_),
    .RESET_B(net287),
    .Q(\line_cache[23][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26552_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00364_),
    .RESET_B(net286),
    .Q(\line_cache[23][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26553_ (.CLK(clknet_leaf_237_clk_i),
    .D(_00365_),
    .RESET_B(net264),
    .Q(\line_cache[23][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26554_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00366_),
    .RESET_B(net286),
    .Q(\line_cache[23][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26555_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00367_),
    .RESET_B(net290),
    .Q(\line_cache[23][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26556_ (.CLK(clknet_leaf_243_clk_i),
    .D(_00368_),
    .RESET_B(net289),
    .Q(\line_cache[23][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26557_ (.CLK(clknet_leaf_240_clk_i),
    .D(_00369_),
    .RESET_B(net287),
    .Q(\line_cache[23][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26558_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00370_),
    .RESET_B(net287),
    .Q(\line_cache[23][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26559_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00371_),
    .RESET_B(net296),
    .Q(\line_cache[24][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26560_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00372_),
    .RESET_B(net292),
    .Q(\line_cache[24][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26561_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00373_),
    .RESET_B(net297),
    .Q(\line_cache[24][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26562_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00374_),
    .RESET_B(net293),
    .Q(\line_cache[24][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26563_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00375_),
    .RESET_B(net297),
    .Q(\line_cache[24][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26564_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00376_),
    .RESET_B(net294),
    .Q(\line_cache[24][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26565_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00377_),
    .RESET_B(net297),
    .Q(\line_cache[24][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26566_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00378_),
    .RESET_B(net292),
    .Q(\line_cache[24][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26567_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00379_),
    .RESET_B(net296),
    .Q(\line_cache[25][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26568_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00380_),
    .RESET_B(net292),
    .Q(\line_cache[25][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26569_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00381_),
    .RESET_B(net296),
    .Q(\line_cache[25][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26570_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00382_),
    .RESET_B(net294),
    .Q(\line_cache[25][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26571_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00383_),
    .RESET_B(net297),
    .Q(\line_cache[25][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26572_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00384_),
    .RESET_B(net294),
    .Q(\line_cache[25][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26573_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00385_),
    .RESET_B(net297),
    .Q(\line_cache[25][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26574_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00386_),
    .RESET_B(net292),
    .Q(\line_cache[25][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26575_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00387_),
    .RESET_B(net296),
    .Q(\line_cache[26][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26576_ (.CLK(clknet_leaf_242_clk_i),
    .D(_00388_),
    .RESET_B(net286),
    .Q(\line_cache[26][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26577_ (.CLK(clknet_leaf_250_clk_i),
    .D(_00389_),
    .RESET_B(net296),
    .Q(\line_cache[26][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26578_ (.CLK(clknet_leaf_256_clk_i),
    .D(_00390_),
    .RESET_B(net294),
    .Q(\line_cache[26][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26579_ (.CLK(clknet_leaf_256_clk_i),
    .D(_00391_),
    .RESET_B(net294),
    .Q(\line_cache[26][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26580_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00392_),
    .RESET_B(net297),
    .Q(\line_cache[26][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26581_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00393_),
    .RESET_B(net297),
    .Q(\line_cache[26][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26582_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00394_),
    .RESET_B(net292),
    .Q(\line_cache[26][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26583_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00395_),
    .RESET_B(net296),
    .Q(\line_cache[27][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26584_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00396_),
    .RESET_B(net292),
    .Q(\line_cache[27][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26585_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00397_),
    .RESET_B(net297),
    .Q(\line_cache[27][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26586_ (.CLK(clknet_leaf_256_clk_i),
    .D(_00398_),
    .RESET_B(net294),
    .Q(\line_cache[27][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26587_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00399_),
    .RESET_B(net297),
    .Q(\line_cache[27][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26588_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00400_),
    .RESET_B(net297),
    .Q(\line_cache[27][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26589_ (.CLK(clknet_leaf_254_clk_i),
    .D(_00401_),
    .RESET_B(net297),
    .Q(\line_cache[27][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26590_ (.CLK(clknet_leaf_255_clk_i),
    .D(_00402_),
    .RESET_B(net296),
    .Q(\line_cache[27][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26591_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00403_),
    .RESET_B(net292),
    .Q(\line_cache[28][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26592_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00404_),
    .RESET_B(net285),
    .Q(\line_cache[28][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26593_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00405_),
    .RESET_B(net295),
    .Q(\line_cache[28][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26594_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00406_),
    .RESET_B(net293),
    .Q(\line_cache[28][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26595_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00407_),
    .RESET_B(net293),
    .Q(\line_cache[28][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26596_ (.CLK(clknet_leaf_256_clk_i),
    .D(_00408_),
    .RESET_B(net294),
    .Q(\line_cache[28][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26597_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00409_),
    .RESET_B(net294),
    .Q(\line_cache[28][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26598_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00410_),
    .RESET_B(net292),
    .Q(\line_cache[28][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26599_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00411_),
    .RESET_B(net295),
    .Q(\line_cache[29][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26600_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00412_),
    .RESET_B(net285),
    .Q(\line_cache[29][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26601_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00413_),
    .RESET_B(net295),
    .Q(\line_cache[29][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26602_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00414_),
    .RESET_B(net293),
    .Q(\line_cache[29][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26603_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00415_),
    .RESET_B(net293),
    .Q(\line_cache[29][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26604_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00416_),
    .RESET_B(net293),
    .Q(\line_cache[29][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26605_ (.CLK(clknet_leaf_256_clk_i),
    .D(_00417_),
    .RESET_B(net294),
    .Q(\line_cache[29][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26606_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00418_),
    .RESET_B(net292),
    .Q(\line_cache[29][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26607_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00419_),
    .RESET_B(net292),
    .Q(\line_cache[30][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26608_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00420_),
    .RESET_B(net292),
    .Q(\line_cache[30][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26609_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00421_),
    .RESET_B(net295),
    .Q(\line_cache[30][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26610_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00422_),
    .RESET_B(net293),
    .Q(\line_cache[30][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26611_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00423_),
    .RESET_B(net293),
    .Q(\line_cache[30][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26612_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00424_),
    .RESET_B(net293),
    .Q(\line_cache[30][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26613_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00425_),
    .RESET_B(net294),
    .Q(\line_cache[30][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26614_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00426_),
    .RESET_B(net292),
    .Q(\line_cache[30][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26615_ (.CLK(clknet_leaf_263_clk_i),
    .D(_00427_),
    .RESET_B(net285),
    .Q(\line_cache[31][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26616_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00428_),
    .RESET_B(net284),
    .Q(\line_cache[31][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26617_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00429_),
    .RESET_B(net284),
    .Q(\line_cache[31][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26618_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00430_),
    .RESET_B(net285),
    .Q(\line_cache[31][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26619_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00431_),
    .RESET_B(net284),
    .Q(\line_cache[31][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26620_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00432_),
    .RESET_B(net285),
    .Q(\line_cache[31][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26621_ (.CLK(clknet_leaf_239_clk_i),
    .D(_00433_),
    .RESET_B(net284),
    .Q(\line_cache[31][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26622_ (.CLK(clknet_leaf_262_clk_i),
    .D(_00434_),
    .RESET_B(net285),
    .Q(\line_cache[31][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26623_ (.CLK(clknet_leaf_261_clk_i),
    .D(_00435_),
    .RESET_B(net295),
    .Q(\line_cache[32][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26624_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00436_),
    .RESET_B(net292),
    .Q(\line_cache[32][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26625_ (.CLK(clknet_leaf_256_clk_i),
    .D(_00437_),
    .RESET_B(net295),
    .Q(\line_cache[32][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26626_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00438_),
    .RESET_B(net293),
    .Q(\line_cache[32][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26627_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00439_),
    .RESET_B(net293),
    .Q(\line_cache[32][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26628_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00440_),
    .RESET_B(net293),
    .Q(\line_cache[32][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26629_ (.CLK(clknet_leaf_257_clk_i),
    .D(_00441_),
    .RESET_B(net294),
    .Q(\line_cache[32][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26630_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00442_),
    .RESET_B(net292),
    .Q(\line_cache[32][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26631_ (.CLK(clknet_leaf_265_clk_i),
    .D(_00443_),
    .RESET_B(net286),
    .Q(\line_cache[33][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26632_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00444_),
    .RESET_B(net280),
    .Q(\line_cache[33][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26633_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00445_),
    .RESET_B(net280),
    .Q(\line_cache[33][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26634_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00446_),
    .RESET_B(net281),
    .Q(\line_cache[33][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26635_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00447_),
    .RESET_B(net281),
    .Q(\line_cache[33][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26636_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00448_),
    .RESET_B(net282),
    .Q(\line_cache[33][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26637_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00449_),
    .RESET_B(net293),
    .Q(\line_cache[33][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26638_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00450_),
    .RESET_B(net280),
    .Q(\line_cache[33][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26639_ (.CLK(clknet_leaf_265_clk_i),
    .D(_00451_),
    .RESET_B(net275),
    .Q(\line_cache[34][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26640_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00452_),
    .RESET_B(net280),
    .Q(\line_cache[34][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26641_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00453_),
    .RESET_B(net280),
    .Q(\line_cache[34][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26642_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00454_),
    .RESET_B(net282),
    .Q(\line_cache[34][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26643_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00455_),
    .RESET_B(net282),
    .Q(\line_cache[34][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26644_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00456_),
    .RESET_B(net282),
    .Q(\line_cache[34][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26645_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00457_),
    .RESET_B(net282),
    .Q(\line_cache[34][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26646_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00458_),
    .RESET_B(net280),
    .Q(\line_cache[34][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26647_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00459_),
    .RESET_B(net280),
    .Q(\line_cache[35][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26648_ (.CLK(clknet_leaf_265_clk_i),
    .D(_00460_),
    .RESET_B(net275),
    .Q(\line_cache[35][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26649_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00461_),
    .RESET_B(net282),
    .Q(\line_cache[35][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26650_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00462_),
    .RESET_B(net282),
    .Q(\line_cache[35][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26651_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00463_),
    .RESET_B(net282),
    .Q(\line_cache[35][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26652_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00464_),
    .RESET_B(net293),
    .Q(\line_cache[35][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26653_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00465_),
    .RESET_B(net293),
    .Q(\line_cache[35][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26654_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00466_),
    .RESET_B(net283),
    .Q(\line_cache[35][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26655_ (.CLK(clknet_leaf_260_clk_i),
    .D(_00467_),
    .RESET_B(net292),
    .Q(\line_cache[36][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26656_ (.CLK(clknet_leaf_265_clk_i),
    .D(_00468_),
    .RESET_B(net275),
    .Q(\line_cache[36][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26657_ (.CLK(clknet_leaf_268_clk_i),
    .D(_00469_),
    .RESET_B(net283),
    .Q(\line_cache[36][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26658_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00470_),
    .RESET_B(net282),
    .Q(\line_cache[36][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26659_ (.CLK(clknet_leaf_269_clk_i),
    .D(_00471_),
    .RESET_B(net282),
    .Q(\line_cache[36][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26660_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00472_),
    .RESET_B(net282),
    .Q(\line_cache[36][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26661_ (.CLK(clknet_leaf_258_clk_i),
    .D(_00473_),
    .RESET_B(net293),
    .Q(\line_cache[36][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26662_ (.CLK(clknet_leaf_259_clk_i),
    .D(_00474_),
    .RESET_B(net292),
    .Q(\line_cache[36][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26663_ (.CLK(clknet_leaf_267_clk_i),
    .D(_00475_),
    .RESET_B(net280),
    .Q(\line_cache[37][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26664_ (.CLK(clknet_leaf_266_clk_i),
    .D(_00476_),
    .RESET_B(net274),
    .Q(\line_cache[37][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26665_ (.CLK(clknet_leaf_267_clk_i),
    .D(_00477_),
    .RESET_B(net280),
    .Q(\line_cache[37][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26666_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00478_),
    .RESET_B(net281),
    .Q(\line_cache[37][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26667_ (.CLK(clknet_leaf_271_clk_i),
    .D(_00479_),
    .RESET_B(net281),
    .Q(\line_cache[37][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26668_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00480_),
    .RESET_B(net279),
    .Q(\line_cache[37][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26669_ (.CLK(clknet_leaf_271_clk_i),
    .D(_00481_),
    .RESET_B(net281),
    .Q(\line_cache[37][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26670_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00482_),
    .RESET_B(net279),
    .Q(\line_cache[37][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26671_ (.CLK(clknet_leaf_267_clk_i),
    .D(_00483_),
    .RESET_B(net280),
    .Q(\line_cache[38][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26672_ (.CLK(clknet_leaf_266_clk_i),
    .D(_00484_),
    .RESET_B(net274),
    .Q(\line_cache[38][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26673_ (.CLK(clknet_leaf_272_clk_i),
    .D(_00485_),
    .RESET_B(net280),
    .Q(\line_cache[38][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26674_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00486_),
    .RESET_B(net281),
    .Q(\line_cache[38][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26675_ (.CLK(clknet_leaf_271_clk_i),
    .D(_00487_),
    .RESET_B(net281),
    .Q(\line_cache[38][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26676_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00488_),
    .RESET_B(net279),
    .Q(\line_cache[38][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26677_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00489_),
    .RESET_B(net279),
    .Q(\line_cache[38][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26678_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00490_),
    .RESET_B(net277),
    .Q(\line_cache[38][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26679_ (.CLK(clknet_leaf_267_clk_i),
    .D(_00491_),
    .RESET_B(net280),
    .Q(\line_cache[39][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26680_ (.CLK(clknet_leaf_266_clk_i),
    .D(_00492_),
    .RESET_B(net274),
    .Q(\line_cache[39][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26681_ (.CLK(clknet_leaf_272_clk_i),
    .D(_00493_),
    .RESET_B(net281),
    .Q(\line_cache[39][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26682_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00494_),
    .RESET_B(net281),
    .Q(\line_cache[39][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26683_ (.CLK(clknet_leaf_271_clk_i),
    .D(_00495_),
    .RESET_B(net281),
    .Q(\line_cache[39][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26684_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00496_),
    .RESET_B(net279),
    .Q(\line_cache[39][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26685_ (.CLK(clknet_leaf_271_clk_i),
    .D(_00497_),
    .RESET_B(net281),
    .Q(\line_cache[39][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26686_ (.CLK(clknet_leaf_272_clk_i),
    .D(_00498_),
    .RESET_B(net280),
    .Q(\line_cache[39][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26687_ (.CLK(clknet_leaf_267_clk_i),
    .D(_00499_),
    .RESET_B(net283),
    .Q(\line_cache[40][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26688_ (.CLK(clknet_leaf_266_clk_i),
    .D(_00500_),
    .RESET_B(net280),
    .Q(\line_cache[40][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26689_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00501_),
    .RESET_B(net281),
    .Q(\line_cache[40][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26690_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00502_),
    .RESET_B(net281),
    .Q(\line_cache[40][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26691_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00503_),
    .RESET_B(net281),
    .Q(\line_cache[40][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26692_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00504_),
    .RESET_B(net279),
    .Q(\line_cache[40][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26693_ (.CLK(clknet_leaf_270_clk_i),
    .D(_00505_),
    .RESET_B(net281),
    .Q(\line_cache[40][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26694_ (.CLK(clknet_leaf_272_clk_i),
    .D(_00506_),
    .RESET_B(net281),
    .Q(\line_cache[40][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26695_ (.CLK(clknet_leaf_278_clk_i),
    .D(_00507_),
    .RESET_B(net277),
    .Q(\line_cache[41][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26696_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00508_),
    .RESET_B(net277),
    .Q(\line_cache[41][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26697_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00509_),
    .RESET_B(net278),
    .Q(\line_cache[41][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26698_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00510_),
    .RESET_B(net279),
    .Q(\line_cache[41][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26699_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00511_),
    .RESET_B(net279),
    .Q(\line_cache[41][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26700_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00512_),
    .RESET_B(net279),
    .Q(\line_cache[41][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26701_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00513_),
    .RESET_B(net278),
    .Q(\line_cache[41][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26702_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00514_),
    .RESET_B(net271),
    .Q(\line_cache[41][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26703_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00515_),
    .RESET_B(net278),
    .Q(\line_cache[42][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26704_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00516_),
    .RESET_B(net277),
    .Q(\line_cache[42][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26705_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00517_),
    .RESET_B(net277),
    .Q(\line_cache[42][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26706_ (.CLK(clknet_leaf_275_clk_i),
    .D(_00518_),
    .RESET_B(net279),
    .Q(\line_cache[42][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26707_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00519_),
    .RESET_B(net279),
    .Q(\line_cache[42][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26708_ (.CLK(clknet_leaf_274_clk_i),
    .D(_00520_),
    .RESET_B(net279),
    .Q(\line_cache[42][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26709_ (.CLK(clknet_leaf_278_clk_i),
    .D(_00521_),
    .RESET_B(net278),
    .Q(\line_cache[42][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26710_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00522_),
    .RESET_B(net278),
    .Q(\line_cache[42][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26711_ (.CLK(clknet_leaf_278_clk_i),
    .D(_00523_),
    .RESET_B(net271),
    .Q(\line_cache[43][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26712_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00524_),
    .RESET_B(net271),
    .Q(\line_cache[43][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26713_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00525_),
    .RESET_B(net277),
    .Q(\line_cache[43][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26714_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00526_),
    .RESET_B(net279),
    .Q(\line_cache[43][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26715_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00527_),
    .RESET_B(net278),
    .Q(\line_cache[43][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26716_ (.CLK(clknet_leaf_273_clk_i),
    .D(_00528_),
    .RESET_B(net278),
    .Q(\line_cache[43][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26717_ (.CLK(clknet_leaf_272_clk_i),
    .D(_00529_),
    .RESET_B(net280),
    .Q(\line_cache[43][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26718_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00530_),
    .RESET_B(net274),
    .Q(\line_cache[43][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26719_ (.CLK(clknet_leaf_278_clk_i),
    .D(_00531_),
    .RESET_B(net271),
    .Q(\line_cache[44][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26720_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00532_),
    .RESET_B(net271),
    .Q(\line_cache[44][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26721_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00533_),
    .RESET_B(net277),
    .Q(\line_cache[44][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26722_ (.CLK(clknet_leaf_276_clk_i),
    .D(_00534_),
    .RESET_B(net277),
    .Q(\line_cache[44][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26723_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00535_),
    .RESET_B(net278),
    .Q(\line_cache[44][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26724_ (.CLK(clknet_leaf_277_clk_i),
    .D(_00536_),
    .RESET_B(net278),
    .Q(\line_cache[44][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26725_ (.CLK(clknet_leaf_267_clk_i),
    .D(_00537_),
    .RESET_B(net280),
    .Q(\line_cache[44][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26726_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00538_),
    .RESET_B(net274),
    .Q(\line_cache[44][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26727_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00539_),
    .RESET_B(net256),
    .Q(\line_cache[45][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26728_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00540_),
    .RESET_B(net256),
    .Q(\line_cache[45][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26729_ (.CLK(clknet_leaf_288_clk_i),
    .D(_00541_),
    .RESET_B(net256),
    .Q(\line_cache[45][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26730_ (.CLK(clknet_leaf_288_clk_i),
    .D(_00542_),
    .RESET_B(net256),
    .Q(\line_cache[45][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26731_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00543_),
    .RESET_B(net273),
    .Q(\line_cache[45][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26732_ (.CLK(clknet_leaf_286_clk_i),
    .D(_00544_),
    .RESET_B(net276),
    .Q(\line_cache[45][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26733_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00545_),
    .RESET_B(net256),
    .Q(\line_cache[45][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26734_ (.CLK(clknet_leaf_286_clk_i),
    .D(_00546_),
    .RESET_B(net276),
    .Q(\line_cache[45][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26735_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00547_),
    .RESET_B(net256),
    .Q(\line_cache[46][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26736_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00548_),
    .RESET_B(net256),
    .Q(\line_cache[46][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26737_ (.CLK(clknet_leaf_288_clk_i),
    .D(_00549_),
    .RESET_B(net256),
    .Q(\line_cache[46][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26738_ (.CLK(clknet_leaf_287_clk_i),
    .D(_00550_),
    .RESET_B(net256),
    .Q(\line_cache[46][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26739_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00551_),
    .RESET_B(net273),
    .Q(\line_cache[46][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26740_ (.CLK(clknet_leaf_286_clk_i),
    .D(_00552_),
    .RESET_B(net276),
    .Q(\line_cache[46][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26741_ (.CLK(clknet_leaf_287_clk_i),
    .D(_00553_),
    .RESET_B(net256),
    .Q(\line_cache[46][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26742_ (.CLK(clknet_leaf_286_clk_i),
    .D(_00554_),
    .RESET_B(net276),
    .Q(\line_cache[46][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26743_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00555_),
    .RESET_B(net264),
    .Q(\line_cache[47][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26744_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00556_),
    .RESET_B(net264),
    .Q(\line_cache[47][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26745_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00557_),
    .RESET_B(net264),
    .Q(\line_cache[47][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26746_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00558_),
    .RESET_B(net264),
    .Q(\line_cache[47][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26747_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00559_),
    .RESET_B(net264),
    .Q(\line_cache[47][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26748_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00560_),
    .RESET_B(net264),
    .Q(\line_cache[47][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26749_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00561_),
    .RESET_B(net268),
    .Q(\line_cache[47][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26750_ (.CLK(clknet_leaf_238_clk_i),
    .D(_00562_),
    .RESET_B(net268),
    .Q(\line_cache[47][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26751_ (.CLK(clknet_leaf_289_clk_i),
    .D(_00563_),
    .RESET_B(net256),
    .Q(\line_cache[48][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26752_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00564_),
    .RESET_B(net253),
    .Q(\line_cache[48][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26753_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00565_),
    .RESET_B(net253),
    .Q(\line_cache[48][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26754_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00566_),
    .RESET_B(net269),
    .Q(\line_cache[48][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26755_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00567_),
    .RESET_B(net269),
    .Q(\line_cache[48][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26756_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00568_),
    .RESET_B(net269),
    .Q(\line_cache[48][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26757_ (.CLK(clknet_leaf_288_clk_i),
    .D(_00569_),
    .RESET_B(net256),
    .Q(\line_cache[48][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26758_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00570_),
    .RESET_B(net273),
    .Q(\line_cache[48][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26759_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00571_),
    .RESET_B(net253),
    .Q(\line_cache[49][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26760_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00572_),
    .RESET_B(net253),
    .Q(\line_cache[49][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26761_ (.CLK(clknet_leaf_293_clk_i),
    .D(_00573_),
    .RESET_B(net254),
    .Q(\line_cache[49][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26762_ (.CLK(clknet_leaf_281_clk_i),
    .D(_00574_),
    .RESET_B(net269),
    .Q(\line_cache[49][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26763_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00575_),
    .RESET_B(net270),
    .Q(\line_cache[49][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26764_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00576_),
    .RESET_B(net270),
    .Q(\line_cache[49][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26765_ (.CLK(clknet_leaf_288_clk_i),
    .D(_00577_),
    .RESET_B(net256),
    .Q(\line_cache[49][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26766_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00578_),
    .RESET_B(net273),
    .Q(\line_cache[49][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26767_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00579_),
    .RESET_B(net254),
    .Q(\line_cache[50][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26768_ (.CLK(clknet_leaf_293_clk_i),
    .D(_00580_),
    .RESET_B(net253),
    .Q(\line_cache[50][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26769_ (.CLK(clknet_leaf_294_clk_i),
    .D(_00581_),
    .RESET_B(net253),
    .Q(\line_cache[50][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26770_ (.CLK(clknet_leaf_281_clk_i),
    .D(_00582_),
    .RESET_B(net269),
    .Q(\line_cache[50][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26771_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00583_),
    .RESET_B(net270),
    .Q(\line_cache[50][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26772_ (.CLK(clknet_leaf_289_clk_i),
    .D(_00584_),
    .RESET_B(net273),
    .Q(\line_cache[50][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26773_ (.CLK(clknet_leaf_289_clk_i),
    .D(_00585_),
    .RESET_B(net256),
    .Q(\line_cache[50][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26774_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00586_),
    .RESET_B(net273),
    .Q(\line_cache[50][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26775_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00587_),
    .RESET_B(net254),
    .Q(\line_cache[51][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26776_ (.CLK(clknet_leaf_293_clk_i),
    .D(_00588_),
    .RESET_B(net253),
    .Q(\line_cache[51][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26777_ (.CLK(clknet_leaf_295_clk_i),
    .D(_00589_),
    .RESET_B(net253),
    .Q(\line_cache[51][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26778_ (.CLK(clknet_leaf_293_clk_i),
    .D(_00590_),
    .RESET_B(net269),
    .Q(\line_cache[51][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26779_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00591_),
    .RESET_B(net270),
    .Q(\line_cache[51][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26780_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00592_),
    .RESET_B(net270),
    .Q(\line_cache[51][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26781_ (.CLK(clknet_leaf_292_clk_i),
    .D(_00593_),
    .RESET_B(net254),
    .Q(\line_cache[51][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26782_ (.CLK(clknet_leaf_284_clk_i),
    .D(_00594_),
    .RESET_B(net273),
    .Q(\line_cache[51][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26783_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00595_),
    .RESET_B(net272),
    .Q(\line_cache[52][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26784_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00596_),
    .RESET_B(net271),
    .Q(\line_cache[52][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26785_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00597_),
    .RESET_B(net272),
    .Q(\line_cache[52][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26786_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00598_),
    .RESET_B(net271),
    .Q(\line_cache[52][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26787_ (.CLK(clknet_leaf_278_clk_i),
    .D(_00599_),
    .RESET_B(net272),
    .Q(\line_cache[52][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26788_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00600_),
    .RESET_B(net274),
    .Q(\line_cache[52][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26789_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00601_),
    .RESET_B(net274),
    .Q(\line_cache[52][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26790_ (.CLK(clknet_leaf_284_clk_i),
    .D(_00602_),
    .RESET_B(net274),
    .Q(\line_cache[52][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26791_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00603_),
    .RESET_B(net272),
    .Q(\line_cache[53][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26792_ (.CLK(clknet_leaf_280_clk_i),
    .D(_00604_),
    .RESET_B(net271),
    .Q(\line_cache[53][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26793_ (.CLK(clknet_leaf_278_clk_i),
    .D(_00605_),
    .RESET_B(net272),
    .Q(\line_cache[53][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26794_ (.CLK(clknet_leaf_279_clk_i),
    .D(_00606_),
    .RESET_B(net271),
    .Q(\line_cache[53][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26795_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00607_),
    .RESET_B(net272),
    .Q(\line_cache[53][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26796_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00608_),
    .RESET_B(net272),
    .Q(\line_cache[53][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26797_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00609_),
    .RESET_B(net274),
    .Q(\line_cache[53][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26798_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00610_),
    .RESET_B(net273),
    .Q(\line_cache[53][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26799_ (.CLK(clknet_leaf_283_clk_i),
    .D(_00611_),
    .RESET_B(net272),
    .Q(\line_cache[54][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26800_ (.CLK(clknet_leaf_281_clk_i),
    .D(_00612_),
    .RESET_B(net269),
    .Q(\line_cache[54][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26801_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00613_),
    .RESET_B(net270),
    .Q(\line_cache[54][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26802_ (.CLK(clknet_leaf_280_clk_i),
    .D(_00614_),
    .RESET_B(net271),
    .Q(\line_cache[54][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26803_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00615_),
    .RESET_B(net272),
    .Q(\line_cache[54][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26804_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00616_),
    .RESET_B(net270),
    .Q(\line_cache[54][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26805_ (.CLK(clknet_leaf_284_clk_i),
    .D(_00617_),
    .RESET_B(net274),
    .Q(\line_cache[54][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26806_ (.CLK(clknet_leaf_285_clk_i),
    .D(_00618_),
    .RESET_B(net273),
    .Q(\line_cache[54][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26807_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00619_),
    .RESET_B(net270),
    .Q(\line_cache[55][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26808_ (.CLK(clknet_leaf_281_clk_i),
    .D(_00620_),
    .RESET_B(net269),
    .Q(\line_cache[55][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26809_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00621_),
    .RESET_B(net269),
    .Q(\line_cache[55][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26810_ (.CLK(clknet_leaf_281_clk_i),
    .D(_00622_),
    .RESET_B(net269),
    .Q(\line_cache[55][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26811_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00623_),
    .RESET_B(net270),
    .Q(\line_cache[55][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26812_ (.CLK(clknet_leaf_282_clk_i),
    .D(_00624_),
    .RESET_B(net270),
    .Q(\line_cache[55][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26813_ (.CLK(clknet_leaf_284_clk_i),
    .D(_00625_),
    .RESET_B(net273),
    .Q(\line_cache[55][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26814_ (.CLK(clknet_leaf_284_clk_i),
    .D(_00626_),
    .RESET_B(net273),
    .Q(\line_cache[55][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26815_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00627_),
    .RESET_B(net254),
    .Q(\line_cache[56][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26816_ (.CLK(clknet_leaf_295_clk_i),
    .D(_00628_),
    .RESET_B(net253),
    .Q(\line_cache[56][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26817_ (.CLK(clknet_leaf_297_clk_i),
    .D(_00629_),
    .RESET_B(net253),
    .Q(\line_cache[56][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26818_ (.CLK(clknet_leaf_295_clk_i),
    .D(_00630_),
    .RESET_B(net251),
    .Q(\line_cache[56][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26819_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00631_),
    .RESET_B(net254),
    .Q(\line_cache[56][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26820_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00632_),
    .RESET_B(net254),
    .Q(\line_cache[56][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26821_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00633_),
    .RESET_B(net256),
    .Q(\line_cache[56][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26822_ (.CLK(clknet_leaf_289_clk_i),
    .D(_00634_),
    .RESET_B(net256),
    .Q(\line_cache[56][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26823_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00635_),
    .RESET_B(net251),
    .Q(\line_cache[57][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26824_ (.CLK(clknet_leaf_295_clk_i),
    .D(_00636_),
    .RESET_B(net251),
    .Q(\line_cache[57][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26825_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00637_),
    .RESET_B(net251),
    .Q(\line_cache[57][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26826_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00638_),
    .RESET_B(net251),
    .Q(\line_cache[57][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26827_ (.CLK(clknet_leaf_291_clk_i),
    .D(_00639_),
    .RESET_B(net252),
    .Q(\line_cache[57][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26828_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00640_),
    .RESET_B(net252),
    .Q(\line_cache[57][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26829_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00641_),
    .RESET_B(net255),
    .Q(\line_cache[57][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26830_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00642_),
    .RESET_B(net255),
    .Q(\line_cache[57][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26831_ (.CLK(clknet_leaf_298_clk_i),
    .D(_00643_),
    .RESET_B(net252),
    .Q(\line_cache[58][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26832_ (.CLK(clknet_leaf_298_clk_i),
    .D(_00644_),
    .RESET_B(net252),
    .Q(\line_cache[58][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26833_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00645_),
    .RESET_B(net251),
    .Q(\line_cache[58][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26834_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00646_),
    .RESET_B(net251),
    .Q(\line_cache[58][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26835_ (.CLK(clknet_leaf_297_clk_i),
    .D(_00647_),
    .RESET_B(net252),
    .Q(\line_cache[58][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26836_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00648_),
    .RESET_B(net252),
    .Q(\line_cache[58][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26837_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00649_),
    .RESET_B(net252),
    .Q(\line_cache[58][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26838_ (.CLK(clknet_leaf_312_clk_i),
    .D(_00650_),
    .RESET_B(net255),
    .Q(\line_cache[58][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26839_ (.CLK(clknet_leaf_306_clk_i),
    .D(_00651_),
    .RESET_B(net252),
    .Q(\line_cache[59][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26840_ (.CLK(clknet_leaf_297_clk_i),
    .D(_00652_),
    .RESET_B(net252),
    .Q(\line_cache[59][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26841_ (.CLK(clknet_leaf_296_clk_i),
    .D(_00653_),
    .RESET_B(net251),
    .Q(\line_cache[59][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26842_ (.CLK(clknet_leaf_298_clk_i),
    .D(_00654_),
    .RESET_B(net252),
    .Q(\line_cache[59][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26843_ (.CLK(clknet_leaf_297_clk_i),
    .D(_00655_),
    .RESET_B(net252),
    .Q(\line_cache[59][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26844_ (.CLK(clknet_leaf_297_clk_i),
    .D(_00656_),
    .RESET_B(net252),
    .Q(\line_cache[59][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26845_ (.CLK(clknet_leaf_290_clk_i),
    .D(_00657_),
    .RESET_B(net255),
    .Q(\line_cache[59][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26846_ (.CLK(clknet_leaf_313_clk_i),
    .D(_00658_),
    .RESET_B(net249),
    .Q(\line_cache[59][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26847_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00659_),
    .RESET_B(net255),
    .Q(\line_cache[60][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26848_ (.CLK(clknet_leaf_313_clk_i),
    .D(_00660_),
    .RESET_B(net255),
    .Q(\line_cache[60][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26849_ (.CLK(clknet_leaf_312_clk_i),
    .D(_00661_),
    .RESET_B(net255),
    .Q(\line_cache[60][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26850_ (.CLK(clknet_leaf_311_clk_i),
    .D(_00662_),
    .RESET_B(net255),
    .Q(\line_cache[60][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26851_ (.CLK(clknet_leaf_313_clk_i),
    .D(_00663_),
    .RESET_B(net255),
    .Q(\line_cache[60][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26852_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00664_),
    .RESET_B(net255),
    .Q(\line_cache[60][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26853_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00665_),
    .RESET_B(net255),
    .Q(\line_cache[60][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26854_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00666_),
    .RESET_B(net257),
    .Q(\line_cache[60][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26855_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00667_),
    .RESET_B(net255),
    .Q(\line_cache[61][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26856_ (.CLK(clknet_leaf_313_clk_i),
    .D(_00668_),
    .RESET_B(net255),
    .Q(\line_cache[61][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26857_ (.CLK(clknet_leaf_312_clk_i),
    .D(_00669_),
    .RESET_B(net255),
    .Q(\line_cache[61][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26858_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00670_),
    .RESET_B(net255),
    .Q(\line_cache[61][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26859_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00671_),
    .RESET_B(net255),
    .Q(\line_cache[61][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26860_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00672_),
    .RESET_B(net257),
    .Q(\line_cache[61][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26861_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00673_),
    .RESET_B(net268),
    .Q(\line_cache[61][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26862_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00674_),
    .RESET_B(net268),
    .Q(\line_cache[61][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26863_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00675_),
    .RESET_B(net257),
    .Q(\line_cache[62][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26864_ (.CLK(clknet_leaf_316_clk_i),
    .D(_00676_),
    .RESET_B(net263),
    .Q(\line_cache[62][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26865_ (.CLK(clknet_leaf_311_clk_i),
    .D(_00677_),
    .RESET_B(net257),
    .Q(\line_cache[62][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26866_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00678_),
    .RESET_B(net257),
    .Q(\line_cache[62][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26867_ (.CLK(clknet_leaf_314_clk_i),
    .D(_00679_),
    .RESET_B(net257),
    .Q(\line_cache[62][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26868_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00680_),
    .RESET_B(net257),
    .Q(\line_cache[62][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26869_ (.CLK(clknet_leaf_316_clk_i),
    .D(_00681_),
    .RESET_B(net263),
    .Q(\line_cache[62][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26870_ (.CLK(clknet_leaf_316_clk_i),
    .D(_00682_),
    .RESET_B(net263),
    .Q(\line_cache[62][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26871_ (.CLK(clknet_leaf_236_clk_i),
    .D(_00683_),
    .RESET_B(net263),
    .Q(\line_cache[63][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26872_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00684_),
    .RESET_B(net263),
    .Q(\line_cache[63][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26873_ (.CLK(clknet_leaf_316_clk_i),
    .D(_00685_),
    .RESET_B(net263),
    .Q(\line_cache[63][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26874_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00686_),
    .RESET_B(net263),
    .Q(\line_cache[63][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26875_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00687_),
    .RESET_B(net264),
    .Q(\line_cache[63][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26876_ (.CLK(clknet_leaf_315_clk_i),
    .D(_00688_),
    .RESET_B(net268),
    .Q(\line_cache[63][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26877_ (.CLK(clknet_leaf_317_clk_i),
    .D(_00689_),
    .RESET_B(net268),
    .Q(\line_cache[63][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26878_ (.CLK(clknet_leaf_316_clk_i),
    .D(_00690_),
    .RESET_B(net263),
    .Q(\line_cache[63][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26879_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00691_),
    .RESET_B(net328),
    .Q(\line_cache[64][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26880_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00692_),
    .RESET_B(net309),
    .Q(\line_cache[64][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26881_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00693_),
    .RESET_B(net328),
    .Q(\line_cache[64][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26882_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00694_),
    .RESET_B(net309),
    .Q(\line_cache[64][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26883_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00695_),
    .RESET_B(net329),
    .Q(\line_cache[64][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26884_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00696_),
    .RESET_B(net309),
    .Q(\line_cache[64][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26885_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00697_),
    .RESET_B(net329),
    .Q(\line_cache[64][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26886_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00698_),
    .RESET_B(net309),
    .Q(\line_cache[64][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26887_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00699_),
    .RESET_B(net328),
    .Q(\line_cache[65][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26888_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00700_),
    .RESET_B(net309),
    .Q(\line_cache[65][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26889_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00701_),
    .RESET_B(net328),
    .Q(\line_cache[65][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26890_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00702_),
    .RESET_B(net309),
    .Q(\line_cache[65][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26891_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00703_),
    .RESET_B(net328),
    .Q(\line_cache[65][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26892_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00704_),
    .RESET_B(net310),
    .Q(\line_cache[65][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26893_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00705_),
    .RESET_B(net328),
    .Q(\line_cache[65][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26894_ (.CLK(clknet_leaf_222_clk_i),
    .D(_00706_),
    .RESET_B(net309),
    .Q(\line_cache[65][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26895_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00707_),
    .RESET_B(net328),
    .Q(\line_cache[66][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26896_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00708_),
    .RESET_B(net310),
    .Q(\line_cache[66][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26897_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00709_),
    .RESET_B(net328),
    .Q(\line_cache[66][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26898_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00710_),
    .RESET_B(net307),
    .Q(\line_cache[66][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26899_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00711_),
    .RESET_B(net329),
    .Q(\line_cache[66][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26900_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00712_),
    .RESET_B(net310),
    .Q(\line_cache[66][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26901_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00713_),
    .RESET_B(net329),
    .Q(\line_cache[66][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26902_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00714_),
    .RESET_B(net309),
    .Q(\line_cache[66][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26903_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00715_),
    .RESET_B(net328),
    .Q(\line_cache[67][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26904_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00716_),
    .RESET_B(net310),
    .Q(\line_cache[67][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26905_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00717_),
    .RESET_B(net328),
    .Q(\line_cache[67][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26906_ (.CLK(clknet_leaf_223_clk_i),
    .D(_00718_),
    .RESET_B(net307),
    .Q(\line_cache[67][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26907_ (.CLK(clknet_leaf_209_clk_i),
    .D(_00719_),
    .RESET_B(net329),
    .Q(\line_cache[67][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26908_ (.CLK(clknet_leaf_224_clk_i),
    .D(_00720_),
    .RESET_B(net309),
    .Q(\line_cache[67][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26909_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00721_),
    .RESET_B(net329),
    .Q(\line_cache[67][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26910_ (.CLK(clknet_leaf_221_clk_i),
    .D(_00722_),
    .RESET_B(net309),
    .Q(\line_cache[67][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26911_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00723_),
    .RESET_B(net333),
    .Q(\line_cache[68][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26912_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00724_),
    .RESET_B(net339),
    .Q(\line_cache[68][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26913_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00725_),
    .RESET_B(net341),
    .Q(\line_cache[68][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26914_ (.CLK(clknet_leaf_194_clk_i),
    .D(_00726_),
    .RESET_B(net339),
    .Q(\line_cache[68][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26915_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00727_),
    .RESET_B(net341),
    .Q(\line_cache[68][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26916_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00728_),
    .RESET_B(net339),
    .Q(\line_cache[68][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26917_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00729_),
    .RESET_B(net341),
    .Q(\line_cache[68][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26918_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00730_),
    .RESET_B(net341),
    .Q(\line_cache[68][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26919_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00731_),
    .RESET_B(net333),
    .Q(\line_cache[69][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26920_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00732_),
    .RESET_B(net339),
    .Q(\line_cache[69][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26921_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00733_),
    .RESET_B(net341),
    .Q(\line_cache[69][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26922_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00734_),
    .RESET_B(net333),
    .Q(\line_cache[69][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26923_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00735_),
    .RESET_B(net341),
    .Q(\line_cache[69][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26924_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00736_),
    .RESET_B(net339),
    .Q(\line_cache[69][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26925_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00737_),
    .RESET_B(net341),
    .Q(\line_cache[69][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26926_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00738_),
    .RESET_B(net341),
    .Q(\line_cache[69][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26927_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00739_),
    .RESET_B(net329),
    .Q(\line_cache[70][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26928_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00740_),
    .RESET_B(net330),
    .Q(\line_cache[70][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26929_ (.CLK(clknet_leaf_194_clk_i),
    .D(_00741_),
    .RESET_B(net339),
    .Q(\line_cache[70][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26930_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00742_),
    .RESET_B(net333),
    .Q(\line_cache[70][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26931_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00743_),
    .RESET_B(net339),
    .Q(\line_cache[70][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26932_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00744_),
    .RESET_B(net333),
    .Q(\line_cache[70][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26933_ (.CLK(clknet_leaf_194_clk_i),
    .D(_00745_),
    .RESET_B(net339),
    .Q(\line_cache[70][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26934_ (.CLK(clknet_leaf_194_clk_i),
    .D(_00746_),
    .RESET_B(net339),
    .Q(\line_cache[70][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26935_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00747_),
    .RESET_B(net330),
    .Q(\line_cache[71][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26936_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00748_),
    .RESET_B(net339),
    .Q(\line_cache[71][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26937_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00749_),
    .RESET_B(net339),
    .Q(\line_cache[71][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26938_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00750_),
    .RESET_B(net333),
    .Q(\line_cache[71][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26939_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00751_),
    .RESET_B(net339),
    .Q(\line_cache[71][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26940_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00752_),
    .RESET_B(net333),
    .Q(\line_cache[71][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26941_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00753_),
    .RESET_B(net339),
    .Q(\line_cache[71][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26942_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00754_),
    .RESET_B(net339),
    .Q(\line_cache[71][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26943_ (.CLK(clknet_leaf_193_clk_i),
    .D(_00755_),
    .RESET_B(net333),
    .Q(\line_cache[72][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26944_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00756_),
    .RESET_B(net313),
    .Q(\line_cache[72][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26945_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00757_),
    .RESET_B(net333),
    .Q(\line_cache[72][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26946_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00758_),
    .RESET_B(net311),
    .Q(\line_cache[72][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26947_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00759_),
    .RESET_B(net333),
    .Q(\line_cache[72][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26948_ (.CLK(clknet_leaf_149_clk_i),
    .D(_00760_),
    .RESET_B(net313),
    .Q(\line_cache[72][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26949_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00761_),
    .RESET_B(net332),
    .Q(\line_cache[72][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26950_ (.CLK(clknet_leaf_152_clk_i),
    .D(_00762_),
    .RESET_B(net332),
    .Q(\line_cache[72][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26951_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00763_),
    .RESET_B(net332),
    .Q(\line_cache[73][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26952_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00764_),
    .RESET_B(net332),
    .Q(\line_cache[73][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26953_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00765_),
    .RESET_B(net332),
    .Q(\line_cache[73][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26954_ (.CLK(clknet_leaf_150_clk_i),
    .D(_00766_),
    .RESET_B(net313),
    .Q(\line_cache[73][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26955_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00767_),
    .RESET_B(net333),
    .Q(\line_cache[73][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26956_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00768_),
    .RESET_B(net313),
    .Q(\line_cache[73][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26957_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00769_),
    .RESET_B(net332),
    .Q(\line_cache[73][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26958_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00770_),
    .RESET_B(net313),
    .Q(\line_cache[73][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26959_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00771_),
    .RESET_B(net334),
    .Q(\line_cache[74][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26960_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00772_),
    .RESET_B(net313),
    .Q(\line_cache[74][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26961_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00773_),
    .RESET_B(net333),
    .Q(\line_cache[74][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26962_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00774_),
    .RESET_B(net314),
    .Q(\line_cache[74][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26963_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00775_),
    .RESET_B(net333),
    .Q(\line_cache[74][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26964_ (.CLK(clknet_leaf_151_clk_i),
    .D(_00776_),
    .RESET_B(net314),
    .Q(\line_cache[74][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26965_ (.CLK(clknet_leaf_191_clk_i),
    .D(_00777_),
    .RESET_B(net334),
    .Q(\line_cache[74][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26966_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00778_),
    .RESET_B(net334),
    .Q(\line_cache[74][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26967_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00779_),
    .RESET_B(net334),
    .Q(\line_cache[75][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26968_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00780_),
    .RESET_B(net314),
    .Q(\line_cache[75][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26969_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00781_),
    .RESET_B(net334),
    .Q(\line_cache[75][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26970_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00782_),
    .RESET_B(net314),
    .Q(\line_cache[75][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26971_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00783_),
    .RESET_B(net332),
    .Q(\line_cache[75][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26972_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00784_),
    .RESET_B(net313),
    .Q(\line_cache[75][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26973_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00785_),
    .RESET_B(net334),
    .Q(\line_cache[75][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26974_ (.CLK(clknet_leaf_215_clk_i),
    .D(_00786_),
    .RESET_B(net334),
    .Q(\line_cache[75][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26975_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00787_),
    .RESET_B(net332),
    .Q(\line_cache[76][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26976_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00788_),
    .RESET_B(net310),
    .Q(\line_cache[76][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26977_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00789_),
    .RESET_B(net333),
    .Q(\line_cache[76][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26978_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00790_),
    .RESET_B(net313),
    .Q(\line_cache[76][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26979_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00791_),
    .RESET_B(net313),
    .Q(\line_cache[76][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26980_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00792_),
    .RESET_B(net311),
    .Q(\line_cache[76][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26981_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00793_),
    .RESET_B(net333),
    .Q(\line_cache[76][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26982_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00794_),
    .RESET_B(net332),
    .Q(\line_cache[76][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26983_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00795_),
    .RESET_B(net332),
    .Q(\line_cache[77][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26984_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00796_),
    .RESET_B(net310),
    .Q(\line_cache[77][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26985_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00797_),
    .RESET_B(net331),
    .Q(\line_cache[77][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26986_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00798_),
    .RESET_B(net313),
    .Q(\line_cache[77][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26987_ (.CLK(clknet_leaf_220_clk_i),
    .D(_00799_),
    .RESET_B(net331),
    .Q(\line_cache[77][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26988_ (.CLK(clknet_leaf_218_clk_i),
    .D(_00800_),
    .RESET_B(net313),
    .Q(\line_cache[77][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26989_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00801_),
    .RESET_B(net332),
    .Q(\line_cache[77][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26990_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00802_),
    .RESET_B(net332),
    .Q(\line_cache[77][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26991_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00803_),
    .RESET_B(net331),
    .Q(\line_cache[78][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26992_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00804_),
    .RESET_B(net310),
    .Q(\line_cache[78][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26993_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00805_),
    .RESET_B(net332),
    .Q(\line_cache[78][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26994_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00806_),
    .RESET_B(net313),
    .Q(\line_cache[78][3] ));
 sky130_fd_sc_hd__dfrtp_1 _26995_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00807_),
    .RESET_B(net332),
    .Q(\line_cache[78][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26996_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00808_),
    .RESET_B(net313),
    .Q(\line_cache[78][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26997_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00809_),
    .RESET_B(net332),
    .Q(\line_cache[78][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26998_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00810_),
    .RESET_B(net313),
    .Q(\line_cache[78][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26999_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00811_),
    .RESET_B(net331),
    .Q(\line_cache[79][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27000_ (.CLK(clknet_leaf_219_clk_i),
    .D(_00812_),
    .RESET_B(net310),
    .Q(\line_cache[79][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27001_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00813_),
    .RESET_B(net330),
    .Q(\line_cache[79][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27002_ (.CLK(clknet_leaf_217_clk_i),
    .D(_00814_),
    .RESET_B(net313),
    .Q(\line_cache[79][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27003_ (.CLK(clknet_leaf_210_clk_i),
    .D(_00815_),
    .RESET_B(net331),
    .Q(\line_cache[79][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27004_ (.CLK(clknet_leaf_216_clk_i),
    .D(_00816_),
    .RESET_B(net313),
    .Q(\line_cache[79][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27005_ (.CLK(clknet_leaf_213_clk_i),
    .D(_00817_),
    .RESET_B(net333),
    .Q(\line_cache[79][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27006_ (.CLK(clknet_leaf_214_clk_i),
    .D(_00818_),
    .RESET_B(net332),
    .Q(\line_cache[79][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27007_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00819_),
    .RESET_B(net330),
    .Q(\line_cache[80][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27008_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00820_),
    .RESET_B(net335),
    .Q(\line_cache[80][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27009_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00821_),
    .RESET_B(net335),
    .Q(\line_cache[80][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27010_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00822_),
    .RESET_B(net341),
    .Q(\line_cache[80][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27011_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00823_),
    .RESET_B(net337),
    .Q(\line_cache[80][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27012_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00824_),
    .RESET_B(net341),
    .Q(\line_cache[80][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27013_ (.CLK(clknet_leaf_198_clk_i),
    .D(_00825_),
    .RESET_B(net341),
    .Q(\line_cache[80][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27014_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00826_),
    .RESET_B(net335),
    .Q(\line_cache[80][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27015_ (.CLK(clknet_leaf_211_clk_i),
    .D(_00827_),
    .RESET_B(net330),
    .Q(\line_cache[81][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27016_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00828_),
    .RESET_B(net330),
    .Q(\line_cache[81][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27017_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00829_),
    .RESET_B(net335),
    .Q(\line_cache[81][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27018_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00830_),
    .RESET_B(net336),
    .Q(\line_cache[81][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27019_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00831_),
    .RESET_B(net337),
    .Q(\line_cache[81][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27020_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00832_),
    .RESET_B(net337),
    .Q(\line_cache[81][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27021_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00833_),
    .RESET_B(net337),
    .Q(\line_cache[81][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27022_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00834_),
    .RESET_B(net336),
    .Q(\line_cache[81][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27023_ (.CLK(clknet_leaf_212_clk_i),
    .D(_00835_),
    .RESET_B(net330),
    .Q(\line_cache[82][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27024_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00836_),
    .RESET_B(net336),
    .Q(\line_cache[82][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27025_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00837_),
    .RESET_B(net336),
    .Q(\line_cache[82][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27026_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00838_),
    .RESET_B(net338),
    .Q(\line_cache[82][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27027_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00839_),
    .RESET_B(net338),
    .Q(\line_cache[82][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27028_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00840_),
    .RESET_B(net338),
    .Q(\line_cache[82][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27029_ (.CLK(clknet_leaf_200_clk_i),
    .D(_00841_),
    .RESET_B(net338),
    .Q(\line_cache[82][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27030_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00842_),
    .RESET_B(net336),
    .Q(\line_cache[82][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27031_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00843_),
    .RESET_B(net330),
    .Q(\line_cache[83][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27032_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00844_),
    .RESET_B(net336),
    .Q(\line_cache[83][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27033_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00845_),
    .RESET_B(net336),
    .Q(\line_cache[83][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27034_ (.CLK(clknet_leaf_199_clk_i),
    .D(_00846_),
    .RESET_B(net336),
    .Q(\line_cache[83][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27035_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00847_),
    .RESET_B(net337),
    .Q(\line_cache[83][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27036_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00848_),
    .RESET_B(net337),
    .Q(\line_cache[83][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27037_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00849_),
    .RESET_B(net338),
    .Q(\line_cache[83][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27038_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00850_),
    .RESET_B(net336),
    .Q(\line_cache[83][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27039_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00851_),
    .RESET_B(net334),
    .Q(\line_cache[84][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27040_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00852_),
    .RESET_B(net339),
    .Q(\line_cache[84][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27041_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00853_),
    .RESET_B(net341),
    .Q(\line_cache[84][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27042_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00854_),
    .RESET_B(net339),
    .Q(\line_cache[84][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27043_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00855_),
    .RESET_B(net341),
    .Q(\line_cache[84][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27044_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00856_),
    .RESET_B(net340),
    .Q(\line_cache[84][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27045_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00857_),
    .RESET_B(net341),
    .Q(\line_cache[84][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27046_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00858_),
    .RESET_B(net340),
    .Q(\line_cache[84][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27047_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00859_),
    .RESET_B(net334),
    .Q(\line_cache[85][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27048_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00860_),
    .RESET_B(net340),
    .Q(\line_cache[85][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27049_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00861_),
    .RESET_B(net341),
    .Q(\line_cache[85][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27050_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00862_),
    .RESET_B(net340),
    .Q(\line_cache[85][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27051_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00863_),
    .RESET_B(net341),
    .Q(\line_cache[85][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27052_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00864_),
    .RESET_B(net340),
    .Q(\line_cache[85][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27053_ (.CLK(clknet_leaf_197_clk_i),
    .D(_00865_),
    .RESET_B(net342),
    .Q(\line_cache[85][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27054_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00866_),
    .RESET_B(net340),
    .Q(\line_cache[85][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27055_ (.CLK(clknet_leaf_192_clk_i),
    .D(_00867_),
    .RESET_B(net334),
    .Q(\line_cache[86][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27056_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00868_),
    .RESET_B(net348),
    .Q(\line_cache[86][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27057_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00869_),
    .RESET_B(net349),
    .Q(\line_cache[86][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27058_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00870_),
    .RESET_B(net348),
    .Q(\line_cache[86][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27059_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00871_),
    .RESET_B(net349),
    .Q(\line_cache[86][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27060_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00872_),
    .RESET_B(net344),
    .Q(\line_cache[86][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27061_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00873_),
    .RESET_B(net349),
    .Q(\line_cache[86][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27062_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00874_),
    .RESET_B(net340),
    .Q(\line_cache[86][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27063_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00875_),
    .RESET_B(net344),
    .Q(\line_cache[87][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27064_ (.CLK(clknet_leaf_195_clk_i),
    .D(_00876_),
    .RESET_B(net340),
    .Q(\line_cache[87][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27065_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00877_),
    .RESET_B(net342),
    .Q(\line_cache[87][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27066_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00878_),
    .RESET_B(net348),
    .Q(\line_cache[87][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27067_ (.CLK(clknet_leaf_196_clk_i),
    .D(_00879_),
    .RESET_B(net342),
    .Q(\line_cache[87][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27068_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00880_),
    .RESET_B(net348),
    .Q(\line_cache[87][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27069_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00881_),
    .RESET_B(net349),
    .Q(\line_cache[87][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27070_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00882_),
    .RESET_B(net348),
    .Q(\line_cache[87][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27071_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00883_),
    .RESET_B(net344),
    .Q(\line_cache[88][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27072_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00884_),
    .RESET_B(net348),
    .Q(\line_cache[88][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27073_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00885_),
    .RESET_B(net349),
    .Q(\line_cache[88][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27074_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00886_),
    .RESET_B(net351),
    .Q(\line_cache[88][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27075_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00887_),
    .RESET_B(net349),
    .Q(\line_cache[88][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27076_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00888_),
    .RESET_B(net351),
    .Q(\line_cache[88][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27077_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00889_),
    .RESET_B(net351),
    .Q(\line_cache[88][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27078_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00890_),
    .RESET_B(net351),
    .Q(\line_cache[88][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27079_ (.CLK(clknet_leaf_175_clk_i),
    .D(_00891_),
    .RESET_B(net344),
    .Q(\line_cache[89][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27080_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00892_),
    .RESET_B(net351),
    .Q(\line_cache[89][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27081_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00893_),
    .RESET_B(net349),
    .Q(\line_cache[89][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27082_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00894_),
    .RESET_B(net351),
    .Q(\line_cache[89][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27083_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00895_),
    .RESET_B(net351),
    .Q(\line_cache[89][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27084_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00896_),
    .RESET_B(net347),
    .Q(\line_cache[89][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27085_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00897_),
    .RESET_B(net351),
    .Q(\line_cache[89][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27086_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00898_),
    .RESET_B(net351),
    .Q(\line_cache[89][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27087_ (.CLK(clknet_leaf_179_clk_i),
    .D(_00899_),
    .RESET_B(net347),
    .Q(\line_cache[90][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27088_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00900_),
    .RESET_B(net348),
    .Q(\line_cache[90][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27089_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00901_),
    .RESET_B(net348),
    .Q(\line_cache[90][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27090_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00902_),
    .RESET_B(net351),
    .Q(\line_cache[90][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27091_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00903_),
    .RESET_B(net352),
    .Q(\line_cache[90][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27092_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00904_),
    .RESET_B(net351),
    .Q(\line_cache[90][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27093_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00905_),
    .RESET_B(net352),
    .Q(\line_cache[90][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27094_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00906_),
    .RESET_B(net351),
    .Q(\line_cache[90][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27095_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00907_),
    .RESET_B(net348),
    .Q(\line_cache[91][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27096_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00908_),
    .RESET_B(net351),
    .Q(\line_cache[91][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27097_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00909_),
    .RESET_B(net349),
    .Q(\line_cache[91][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27098_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00910_),
    .RESET_B(net351),
    .Q(\line_cache[91][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27099_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00911_),
    .RESET_B(net349),
    .Q(\line_cache[91][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27100_ (.CLK(clknet_leaf_180_clk_i),
    .D(_00912_),
    .RESET_B(net351),
    .Q(\line_cache[91][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27101_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00913_),
    .RESET_B(net352),
    .Q(\line_cache[91][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27102_ (.CLK(clknet_leaf_181_clk_i),
    .D(_00914_),
    .RESET_B(net351),
    .Q(\line_cache[91][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27103_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00915_),
    .RESET_B(net344),
    .Q(\line_cache[92][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27104_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00916_),
    .RESET_B(net348),
    .Q(\line_cache[92][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27105_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00917_),
    .RESET_B(net349),
    .Q(\line_cache[92][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27106_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00918_),
    .RESET_B(net350),
    .Q(\line_cache[92][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27107_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00919_),
    .RESET_B(net349),
    .Q(\line_cache[92][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27108_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00920_),
    .RESET_B(net350),
    .Q(\line_cache[92][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27109_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00921_),
    .RESET_B(net350),
    .Q(\line_cache[92][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27110_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00922_),
    .RESET_B(net350),
    .Q(\line_cache[92][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27111_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00923_),
    .RESET_B(net350),
    .Q(\line_cache[93][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27112_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00924_),
    .RESET_B(net350),
    .Q(\line_cache[93][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27113_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00925_),
    .RESET_B(net348),
    .Q(\line_cache[93][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27114_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00926_),
    .RESET_B(net348),
    .Q(\line_cache[93][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27115_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00927_),
    .RESET_B(net349),
    .Q(\line_cache[93][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27116_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00928_),
    .RESET_B(net348),
    .Q(\line_cache[93][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27117_ (.CLK(clknet_leaf_183_clk_i),
    .D(_00929_),
    .RESET_B(net350),
    .Q(\line_cache[93][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27118_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00930_),
    .RESET_B(net350),
    .Q(\line_cache[93][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27119_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00931_),
    .RESET_B(net344),
    .Q(\line_cache[94][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27120_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00932_),
    .RESET_B(net350),
    .Q(\line_cache[94][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27121_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00933_),
    .RESET_B(net349),
    .Q(\line_cache[94][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27122_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00934_),
    .RESET_B(net348),
    .Q(\line_cache[94][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27123_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00935_),
    .RESET_B(net349),
    .Q(\line_cache[94][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27124_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00936_),
    .RESET_B(net344),
    .Q(\line_cache[94][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27125_ (.CLK(clknet_leaf_184_clk_i),
    .D(_00937_),
    .RESET_B(net350),
    .Q(\line_cache[94][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27126_ (.CLK(clknet_leaf_182_clk_i),
    .D(_00938_),
    .RESET_B(net350),
    .Q(\line_cache[94][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27127_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00939_),
    .RESET_B(net344),
    .Q(\line_cache[95][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27128_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00940_),
    .RESET_B(net350),
    .Q(\line_cache[95][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27129_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00941_),
    .RESET_B(net349),
    .Q(\line_cache[95][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27130_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00942_),
    .RESET_B(net348),
    .Q(\line_cache[95][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27131_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00943_),
    .RESET_B(net349),
    .Q(\line_cache[95][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27132_ (.CLK(clknet_leaf_186_clk_i),
    .D(_00944_),
    .RESET_B(net348),
    .Q(\line_cache[95][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27133_ (.CLK(clknet_leaf_185_clk_i),
    .D(_00945_),
    .RESET_B(net350),
    .Q(\line_cache[95][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27134_ (.CLK(clknet_leaf_187_clk_i),
    .D(_00946_),
    .RESET_B(net350),
    .Q(\line_cache[95][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27135_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00947_),
    .RESET_B(net330),
    .Q(\line_cache[96][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27136_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00948_),
    .RESET_B(net336),
    .Q(\line_cache[96][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27137_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00949_),
    .RESET_B(net338),
    .Q(\line_cache[96][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27138_ (.CLK(clknet_leaf_205_clk_i),
    .D(_00950_),
    .RESET_B(net335),
    .Q(\line_cache[96][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27139_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00951_),
    .RESET_B(net337),
    .Q(\line_cache[96][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27140_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00952_),
    .RESET_B(net330),
    .Q(\line_cache[96][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27141_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00953_),
    .RESET_B(net337),
    .Q(\line_cache[96][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27142_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00954_),
    .RESET_B(net335),
    .Q(\line_cache[96][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27143_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00955_),
    .RESET_B(net329),
    .Q(\line_cache[97][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27144_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00956_),
    .RESET_B(net335),
    .Q(\line_cache[97][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27145_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00957_),
    .RESET_B(net337),
    .Q(\line_cache[97][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27146_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00958_),
    .RESET_B(net335),
    .Q(\line_cache[97][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27147_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00959_),
    .RESET_B(net337),
    .Q(\line_cache[97][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27148_ (.CLK(clknet_leaf_206_clk_i),
    .D(_00960_),
    .RESET_B(net330),
    .Q(\line_cache[97][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27149_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00961_),
    .RESET_B(net337),
    .Q(\line_cache[97][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27150_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00962_),
    .RESET_B(net335),
    .Q(\line_cache[97][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27151_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00963_),
    .RESET_B(net329),
    .Q(\line_cache[98][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27152_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00964_),
    .RESET_B(net335),
    .Q(\line_cache[98][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27153_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00965_),
    .RESET_B(net337),
    .Q(\line_cache[98][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27154_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00966_),
    .RESET_B(net335),
    .Q(\line_cache[98][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27155_ (.CLK(clknet_leaf_253_clk_i),
    .D(_00967_),
    .RESET_B(net298),
    .Q(\line_cache[98][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27156_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00968_),
    .RESET_B(net329),
    .Q(\line_cache[98][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27157_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00969_),
    .RESET_B(net298),
    .Q(\line_cache[98][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27158_ (.CLK(clknet_leaf_204_clk_i),
    .D(_00970_),
    .RESET_B(net335),
    .Q(\line_cache[98][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27159_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00971_),
    .RESET_B(net329),
    .Q(\line_cache[99][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27160_ (.CLK(clknet_leaf_207_clk_i),
    .D(_00972_),
    .RESET_B(net335),
    .Q(\line_cache[99][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27161_ (.CLK(clknet_leaf_201_clk_i),
    .D(_00973_),
    .RESET_B(net337),
    .Q(\line_cache[99][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27162_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00974_),
    .RESET_B(net337),
    .Q(\line_cache[99][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27163_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00975_),
    .RESET_B(net337),
    .Q(\line_cache[99][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27164_ (.CLK(clknet_leaf_208_clk_i),
    .D(_00976_),
    .RESET_B(net329),
    .Q(\line_cache[99][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27165_ (.CLK(clknet_leaf_202_clk_i),
    .D(_00977_),
    .RESET_B(net337),
    .Q(\line_cache[99][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27166_ (.CLK(clknet_leaf_203_clk_i),
    .D(_00978_),
    .RESET_B(net335),
    .Q(\line_cache[99][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27167_ (.CLK(clknet_leaf_188_clk_i),
    .D(_00979_),
    .RESET_B(net345),
    .Q(\line_cache[100][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27168_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00980_),
    .RESET_B(net334),
    .Q(\line_cache[100][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27169_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00981_),
    .RESET_B(net343),
    .Q(\line_cache[100][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27170_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00982_),
    .RESET_B(net343),
    .Q(\line_cache[100][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27171_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00983_),
    .RESET_B(net344),
    .Q(\line_cache[100][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27172_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00984_),
    .RESET_B(net343),
    .Q(\line_cache[100][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27173_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00985_),
    .RESET_B(net344),
    .Q(\line_cache[100][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27174_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00986_),
    .RESET_B(net343),
    .Q(\line_cache[100][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27175_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00987_),
    .RESET_B(net345),
    .Q(\line_cache[101][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27176_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00988_),
    .RESET_B(net344),
    .Q(\line_cache[101][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27177_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00989_),
    .RESET_B(net343),
    .Q(\line_cache[101][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27178_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00990_),
    .RESET_B(net343),
    .Q(\line_cache[101][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27179_ (.CLK(clknet_leaf_189_clk_i),
    .D(_00991_),
    .RESET_B(net344),
    .Q(\line_cache[101][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27180_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00992_),
    .RESET_B(net343),
    .Q(\line_cache[101][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27181_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00993_),
    .RESET_B(net344),
    .Q(\line_cache[101][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27182_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00994_),
    .RESET_B(net343),
    .Q(\line_cache[101][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27183_ (.CLK(clknet_leaf_174_clk_i),
    .D(_00995_),
    .RESET_B(net343),
    .Q(\line_cache[102][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27184_ (.CLK(clknet_leaf_190_clk_i),
    .D(_00996_),
    .RESET_B(net344),
    .Q(\line_cache[102][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27185_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00997_),
    .RESET_B(net343),
    .Q(\line_cache[102][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27186_ (.CLK(clknet_leaf_172_clk_i),
    .D(_00998_),
    .RESET_B(net343),
    .Q(\line_cache[102][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27187_ (.CLK(clknet_leaf_173_clk_i),
    .D(_00999_),
    .RESET_B(net343),
    .Q(\line_cache[102][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27188_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01000_),
    .RESET_B(net345),
    .Q(\line_cache[102][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27189_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01001_),
    .RESET_B(net343),
    .Q(\line_cache[102][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27190_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01002_),
    .RESET_B(net345),
    .Q(\line_cache[102][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27191_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01003_),
    .RESET_B(net345),
    .Q(\line_cache[103][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27192_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01004_),
    .RESET_B(net344),
    .Q(\line_cache[103][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27193_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01005_),
    .RESET_B(net343),
    .Q(\line_cache[103][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27194_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01006_),
    .RESET_B(net343),
    .Q(\line_cache[103][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27195_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01007_),
    .RESET_B(net345),
    .Q(\line_cache[103][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27196_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01008_),
    .RESET_B(net343),
    .Q(\line_cache[103][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27197_ (.CLK(clknet_leaf_190_clk_i),
    .D(_01009_),
    .RESET_B(net344),
    .Q(\line_cache[103][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27198_ (.CLK(clknet_leaf_173_clk_i),
    .D(_01010_),
    .RESET_B(net345),
    .Q(\line_cache[103][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27199_ (.CLK(clknet_leaf_170_clk_i),
    .D(_01011_),
    .RESET_B(net322),
    .Q(\line_cache[104][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27200_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01012_),
    .RESET_B(net326),
    .Q(\line_cache[104][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27201_ (.CLK(clknet_leaf_170_clk_i),
    .D(_01013_),
    .RESET_B(net324),
    .Q(\line_cache[104][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27202_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01014_),
    .RESET_B(net326),
    .Q(\line_cache[104][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27203_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01015_),
    .RESET_B(net327),
    .Q(\line_cache[104][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27204_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01016_),
    .RESET_B(net326),
    .Q(\line_cache[104][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27205_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01017_),
    .RESET_B(net326),
    .Q(\line_cache[104][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27206_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01018_),
    .RESET_B(net326),
    .Q(\line_cache[104][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27207_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01019_),
    .RESET_B(net324),
    .Q(\line_cache[105][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27208_ (.CLK(clknet_leaf_168_clk_i),
    .D(_01020_),
    .RESET_B(net346),
    .Q(\line_cache[105][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27209_ (.CLK(clknet_leaf_177_clk_i),
    .D(_01021_),
    .RESET_B(net346),
    .Q(\line_cache[105][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27210_ (.CLK(clknet_leaf_168_clk_i),
    .D(_01022_),
    .RESET_B(net327),
    .Q(\line_cache[105][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27211_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01023_),
    .RESET_B(net327),
    .Q(\line_cache[105][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27212_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01024_),
    .RESET_B(net346),
    .Q(\line_cache[105][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27213_ (.CLK(clknet_leaf_177_clk_i),
    .D(_01025_),
    .RESET_B(net346),
    .Q(\line_cache[105][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27214_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01026_),
    .RESET_B(net327),
    .Q(\line_cache[105][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27215_ (.CLK(clknet_leaf_168_clk_i),
    .D(_01027_),
    .RESET_B(net324),
    .Q(\line_cache[106][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27216_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01028_),
    .RESET_B(net346),
    .Q(\line_cache[106][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27217_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01029_),
    .RESET_B(net324),
    .Q(\line_cache[106][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27218_ (.CLK(clknet_leaf_168_clk_i),
    .D(_01030_),
    .RESET_B(net327),
    .Q(\line_cache[106][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27219_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01031_),
    .RESET_B(net327),
    .Q(\line_cache[106][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27220_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01032_),
    .RESET_B(net327),
    .Q(\line_cache[106][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27221_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01033_),
    .RESET_B(net327),
    .Q(\line_cache[106][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27222_ (.CLK(clknet_leaf_168_clk_i),
    .D(_01034_),
    .RESET_B(net327),
    .Q(\line_cache[106][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27223_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01035_),
    .RESET_B(net324),
    .Q(\line_cache[107][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27224_ (.CLK(clknet_leaf_168_clk_i),
    .D(_01036_),
    .RESET_B(net327),
    .Q(\line_cache[107][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27225_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01037_),
    .RESET_B(net324),
    .Q(\line_cache[107][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27226_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01038_),
    .RESET_B(net327),
    .Q(\line_cache[107][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27227_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01039_),
    .RESET_B(net327),
    .Q(\line_cache[107][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27228_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01040_),
    .RESET_B(net353),
    .Q(\line_cache[107][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27229_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01041_),
    .RESET_B(net346),
    .Q(\line_cache[107][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27230_ (.CLK(clknet_leaf_167_clk_i),
    .D(_01042_),
    .RESET_B(net353),
    .Q(\line_cache[107][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27231_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01043_),
    .RESET_B(net345),
    .Q(\line_cache[108][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27232_ (.CLK(clknet_leaf_175_clk_i),
    .D(_01044_),
    .RESET_B(net347),
    .Q(\line_cache[108][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27233_ (.CLK(clknet_leaf_173_clk_i),
    .D(_01045_),
    .RESET_B(net345),
    .Q(\line_cache[108][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27234_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01046_),
    .RESET_B(net347),
    .Q(\line_cache[108][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27235_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01047_),
    .RESET_B(net347),
    .Q(\line_cache[108][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27236_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01048_),
    .RESET_B(net346),
    .Q(\line_cache[108][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27237_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01049_),
    .RESET_B(net347),
    .Q(\line_cache[108][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27238_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01050_),
    .RESET_B(net347),
    .Q(\line_cache[108][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27239_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01051_),
    .RESET_B(net345),
    .Q(\line_cache[109][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27240_ (.CLK(clknet_leaf_176_clk_i),
    .D(_01052_),
    .RESET_B(net347),
    .Q(\line_cache[109][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27241_ (.CLK(clknet_leaf_173_clk_i),
    .D(_01053_),
    .RESET_B(net345),
    .Q(\line_cache[109][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27242_ (.CLK(clknet_leaf_177_clk_i),
    .D(_01054_),
    .RESET_B(net346),
    .Q(\line_cache[109][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27243_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01055_),
    .RESET_B(net347),
    .Q(\line_cache[109][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27244_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01056_),
    .RESET_B(net346),
    .Q(\line_cache[109][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27245_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01057_),
    .RESET_B(net347),
    .Q(\line_cache[109][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27246_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01058_),
    .RESET_B(net346),
    .Q(\line_cache[109][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27247_ (.CLK(clknet_leaf_175_clk_i),
    .D(_01059_),
    .RESET_B(net347),
    .Q(\line_cache[110][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27248_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01060_),
    .RESET_B(net347),
    .Q(\line_cache[110][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27249_ (.CLK(clknet_leaf_173_clk_i),
    .D(_01061_),
    .RESET_B(net345),
    .Q(\line_cache[110][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27250_ (.CLK(clknet_leaf_177_clk_i),
    .D(_01062_),
    .RESET_B(net346),
    .Q(\line_cache[110][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27251_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01063_),
    .RESET_B(net347),
    .Q(\line_cache[110][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27252_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01064_),
    .RESET_B(net352),
    .Q(\line_cache[110][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27253_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01065_),
    .RESET_B(net347),
    .Q(\line_cache[110][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27254_ (.CLK(clknet_leaf_176_clk_i),
    .D(_01066_),
    .RESET_B(net346),
    .Q(\line_cache[110][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27255_ (.CLK(clknet_leaf_174_clk_i),
    .D(_01067_),
    .RESET_B(net345),
    .Q(\line_cache[111][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27256_ (.CLK(clknet_leaf_175_clk_i),
    .D(_01068_),
    .RESET_B(net347),
    .Q(\line_cache[111][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27257_ (.CLK(clknet_leaf_176_clk_i),
    .D(_01069_),
    .RESET_B(net346),
    .Q(\line_cache[111][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27258_ (.CLK(clknet_leaf_176_clk_i),
    .D(_01070_),
    .RESET_B(net346),
    .Q(\line_cache[111][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27259_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01071_),
    .RESET_B(net352),
    .Q(\line_cache[111][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27260_ (.CLK(clknet_leaf_177_clk_i),
    .D(_01072_),
    .RESET_B(net346),
    .Q(\line_cache[111][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27261_ (.CLK(clknet_leaf_179_clk_i),
    .D(_01073_),
    .RESET_B(net347),
    .Q(\line_cache[111][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27262_ (.CLK(clknet_leaf_178_clk_i),
    .D(_01074_),
    .RESET_B(net346),
    .Q(\line_cache[111][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27263_ (.CLK(clknet_leaf_218_clk_i),
    .D(_01075_),
    .RESET_B(net311),
    .Q(\line_cache[112][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27264_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01076_),
    .RESET_B(net307),
    .Q(\line_cache[112][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27265_ (.CLK(clknet_leaf_218_clk_i),
    .D(_01077_),
    .RESET_B(net307),
    .Q(\line_cache[112][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27266_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01078_),
    .RESET_B(net307),
    .Q(\line_cache[112][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27267_ (.CLK(clknet_leaf_219_clk_i),
    .D(_01079_),
    .RESET_B(net308),
    .Q(\line_cache[112][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27268_ (.CLK(clknet_leaf_219_clk_i),
    .D(_01080_),
    .RESET_B(net308),
    .Q(\line_cache[112][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27269_ (.CLK(clknet_leaf_219_clk_i),
    .D(_01081_),
    .RESET_B(net308),
    .Q(\line_cache[112][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27270_ (.CLK(clknet_leaf_218_clk_i),
    .D(_01082_),
    .RESET_B(net311),
    .Q(\line_cache[112][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27271_ (.CLK(clknet_leaf_218_clk_i),
    .D(_01083_),
    .RESET_B(net311),
    .Q(\line_cache[113][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27272_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01084_),
    .RESET_B(net308),
    .Q(\line_cache[113][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27273_ (.CLK(clknet_leaf_218_clk_i),
    .D(_01085_),
    .RESET_B(net308),
    .Q(\line_cache[113][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27274_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01086_),
    .RESET_B(net307),
    .Q(\line_cache[113][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27275_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01087_),
    .RESET_B(net307),
    .Q(\line_cache[113][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27276_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01088_),
    .RESET_B(net308),
    .Q(\line_cache[113][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27277_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01089_),
    .RESET_B(net308),
    .Q(\line_cache[113][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27278_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01090_),
    .RESET_B(net311),
    .Q(\line_cache[113][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27279_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01091_),
    .RESET_B(net311),
    .Q(\line_cache[114][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27280_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01092_),
    .RESET_B(net307),
    .Q(\line_cache[114][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27281_ (.CLK(clknet_leaf_143_clk_i),
    .D(_01093_),
    .RESET_B(net302),
    .Q(\line_cache[114][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27282_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01094_),
    .RESET_B(net302),
    .Q(\line_cache[114][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27283_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01095_),
    .RESET_B(net308),
    .Q(\line_cache[114][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27284_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01096_),
    .RESET_B(net302),
    .Q(\line_cache[114][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27285_ (.CLK(clknet_leaf_143_clk_i),
    .D(_01097_),
    .RESET_B(net302),
    .Q(\line_cache[114][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27286_ (.CLK(clknet_leaf_144_clk_i),
    .D(_01098_),
    .RESET_B(net306),
    .Q(\line_cache[114][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27287_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01099_),
    .RESET_B(net306),
    .Q(\line_cache[115][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27288_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01100_),
    .RESET_B(net308),
    .Q(\line_cache[115][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27289_ (.CLK(clknet_leaf_143_clk_i),
    .D(_01101_),
    .RESET_B(net306),
    .Q(\line_cache[115][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27290_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01102_),
    .RESET_B(net302),
    .Q(\line_cache[115][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27291_ (.CLK(clknet_leaf_225_clk_i),
    .D(_01103_),
    .RESET_B(net308),
    .Q(\line_cache[115][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27292_ (.CLK(clknet_leaf_224_clk_i),
    .D(_01104_),
    .RESET_B(net308),
    .Q(\line_cache[115][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27293_ (.CLK(clknet_leaf_143_clk_i),
    .D(_01105_),
    .RESET_B(net303),
    .Q(\line_cache[115][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27294_ (.CLK(clknet_leaf_144_clk_i),
    .D(_01106_),
    .RESET_B(net306),
    .Q(\line_cache[115][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27295_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01107_),
    .RESET_B(net311),
    .Q(\line_cache[116][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27296_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01108_),
    .RESET_B(net311),
    .Q(\line_cache[116][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27297_ (.CLK(clknet_leaf_144_clk_i),
    .D(_01109_),
    .RESET_B(net306),
    .Q(\line_cache[116][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27298_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01110_),
    .RESET_B(net306),
    .Q(\line_cache[116][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27299_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01111_),
    .RESET_B(net311),
    .Q(\line_cache[116][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27300_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01112_),
    .RESET_B(net311),
    .Q(\line_cache[116][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27301_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01113_),
    .RESET_B(net311),
    .Q(\line_cache[116][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27302_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01114_),
    .RESET_B(net311),
    .Q(\line_cache[116][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27303_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01115_),
    .RESET_B(net312),
    .Q(\line_cache[117][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27304_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01116_),
    .RESET_B(net312),
    .Q(\line_cache[117][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27305_ (.CLK(clknet_leaf_144_clk_i),
    .D(_01117_),
    .RESET_B(net306),
    .Q(\line_cache[117][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27306_ (.CLK(clknet_leaf_144_clk_i),
    .D(_01118_),
    .RESET_B(net306),
    .Q(\line_cache[117][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27307_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01119_),
    .RESET_B(net312),
    .Q(\line_cache[117][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27308_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01120_),
    .RESET_B(net311),
    .Q(\line_cache[117][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27309_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01121_),
    .RESET_B(net306),
    .Q(\line_cache[117][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27310_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01122_),
    .RESET_B(net306),
    .Q(\line_cache[117][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27311_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01123_),
    .RESET_B(net306),
    .Q(\line_cache[118][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27312_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01124_),
    .RESET_B(net312),
    .Q(\line_cache[118][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27313_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01125_),
    .RESET_B(net306),
    .Q(\line_cache[118][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27314_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01126_),
    .RESET_B(net306),
    .Q(\line_cache[118][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27315_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01127_),
    .RESET_B(net312),
    .Q(\line_cache[118][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27316_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01128_),
    .RESET_B(net311),
    .Q(\line_cache[118][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27317_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01129_),
    .RESET_B(net304),
    .Q(\line_cache[118][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27318_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01130_),
    .RESET_B(net306),
    .Q(\line_cache[118][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27319_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01131_),
    .RESET_B(net312),
    .Q(\line_cache[119][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27320_ (.CLK(clknet_leaf_149_clk_i),
    .D(_01132_),
    .RESET_B(net312),
    .Q(\line_cache[119][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27321_ (.CLK(clknet_leaf_145_clk_i),
    .D(_01133_),
    .RESET_B(net304),
    .Q(\line_cache[119][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27322_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01134_),
    .RESET_B(net306),
    .Q(\line_cache[119][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27323_ (.CLK(clknet_leaf_147_clk_i),
    .D(_01135_),
    .RESET_B(net312),
    .Q(\line_cache[119][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27324_ (.CLK(clknet_leaf_148_clk_i),
    .D(_01136_),
    .RESET_B(net311),
    .Q(\line_cache[119][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27325_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01137_),
    .RESET_B(net306),
    .Q(\line_cache[119][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27326_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01138_),
    .RESET_B(net304),
    .Q(\line_cache[119][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27327_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01139_),
    .RESET_B(net322),
    .Q(\line_cache[120][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27328_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01140_),
    .RESET_B(net322),
    .Q(\line_cache[120][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27329_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01141_),
    .RESET_B(net317),
    .Q(\line_cache[120][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27330_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01142_),
    .RESET_B(net315),
    .Q(\line_cache[120][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27331_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01143_),
    .RESET_B(net322),
    .Q(\line_cache[120][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27332_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01144_),
    .RESET_B(net312),
    .Q(\line_cache[120][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27333_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01145_),
    .RESET_B(net323),
    .Q(\line_cache[120][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27334_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01146_),
    .RESET_B(net323),
    .Q(\line_cache[120][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27335_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01147_),
    .RESET_B(net317),
    .Q(\line_cache[121][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27336_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01148_),
    .RESET_B(net323),
    .Q(\line_cache[121][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27337_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01149_),
    .RESET_B(net317),
    .Q(\line_cache[121][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27338_ (.CLK(clknet_leaf_146_clk_i),
    .D(_01150_),
    .RESET_B(net315),
    .Q(\line_cache[121][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27339_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01151_),
    .RESET_B(net322),
    .Q(\line_cache[121][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27340_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01152_),
    .RESET_B(net322),
    .Q(\line_cache[121][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27341_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01153_),
    .RESET_B(net317),
    .Q(\line_cache[121][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27342_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01154_),
    .RESET_B(net317),
    .Q(\line_cache[121][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27343_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01155_),
    .RESET_B(net317),
    .Q(\line_cache[122][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27344_ (.CLK(clknet_leaf_155_clk_i),
    .D(_01156_),
    .RESET_B(net322),
    .Q(\line_cache[122][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27345_ (.CLK(clknet_leaf_155_clk_i),
    .D(_01157_),
    .RESET_B(net317),
    .Q(\line_cache[122][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27346_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01158_),
    .RESET_B(net305),
    .Q(\line_cache[122][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27347_ (.CLK(clknet_leaf_155_clk_i),
    .D(_01159_),
    .RESET_B(net317),
    .Q(\line_cache[122][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27348_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01160_),
    .RESET_B(net322),
    .Q(\line_cache[122][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27349_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01161_),
    .RESET_B(net317),
    .Q(\line_cache[122][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27350_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01162_),
    .RESET_B(net317),
    .Q(\line_cache[122][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27351_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01163_),
    .RESET_B(net323),
    .Q(\line_cache[123][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27352_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01164_),
    .RESET_B(net322),
    .Q(\line_cache[123][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27353_ (.CLK(clknet_leaf_155_clk_i),
    .D(_01165_),
    .RESET_B(net317),
    .Q(\line_cache[123][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27354_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01166_),
    .RESET_B(net317),
    .Q(\line_cache[123][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27355_ (.CLK(clknet_leaf_155_clk_i),
    .D(_01167_),
    .RESET_B(net322),
    .Q(\line_cache[123][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27356_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01168_),
    .RESET_B(net317),
    .Q(\line_cache[123][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27357_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01169_),
    .RESET_B(net317),
    .Q(\line_cache[123][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27358_ (.CLK(clknet_leaf_155_clk_i),
    .D(_01170_),
    .RESET_B(net317),
    .Q(\line_cache[123][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27359_ (.CLK(clknet_leaf_173_clk_i),
    .D(_01171_),
    .RESET_B(net325),
    .Q(\line_cache[124][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27360_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01172_),
    .RESET_B(net324),
    .Q(\line_cache[124][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27361_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01173_),
    .RESET_B(net325),
    .Q(\line_cache[124][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27362_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01174_),
    .RESET_B(net314),
    .Q(\line_cache[124][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27363_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01175_),
    .RESET_B(net324),
    .Q(\line_cache[124][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27364_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01176_),
    .RESET_B(net324),
    .Q(\line_cache[124][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27365_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01177_),
    .RESET_B(net324),
    .Q(\line_cache[124][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27366_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01178_),
    .RESET_B(net325),
    .Q(\line_cache[124][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27367_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01179_),
    .RESET_B(net325),
    .Q(\line_cache[125][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27368_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01180_),
    .RESET_B(net324),
    .Q(\line_cache[125][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27369_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01181_),
    .RESET_B(net325),
    .Q(\line_cache[125][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27370_ (.CLK(clknet_leaf_151_clk_i),
    .D(_01182_),
    .RESET_B(net314),
    .Q(\line_cache[125][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27371_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01183_),
    .RESET_B(net324),
    .Q(\line_cache[125][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27372_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01184_),
    .RESET_B(net324),
    .Q(\line_cache[125][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27373_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01185_),
    .RESET_B(net324),
    .Q(\line_cache[125][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27374_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01186_),
    .RESET_B(net325),
    .Q(\line_cache[125][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27375_ (.CLK(clknet_leaf_170_clk_i),
    .D(_01187_),
    .RESET_B(net323),
    .Q(\line_cache[126][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27376_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01188_),
    .RESET_B(net322),
    .Q(\line_cache[126][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27377_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01189_),
    .RESET_B(net323),
    .Q(\line_cache[126][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27378_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01190_),
    .RESET_B(net312),
    .Q(\line_cache[126][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27379_ (.CLK(clknet_leaf_152_clk_i),
    .D(_01191_),
    .RESET_B(net324),
    .Q(\line_cache[126][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27380_ (.CLK(clknet_leaf_151_clk_i),
    .D(_01192_),
    .RESET_B(net314),
    .Q(\line_cache[126][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27381_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01193_),
    .RESET_B(net322),
    .Q(\line_cache[126][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27382_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01194_),
    .RESET_B(net323),
    .Q(\line_cache[126][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27383_ (.CLK(clknet_leaf_171_clk_i),
    .D(_01195_),
    .RESET_B(net325),
    .Q(\line_cache[127][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27384_ (.CLK(clknet_leaf_172_clk_i),
    .D(_01196_),
    .RESET_B(net324),
    .Q(\line_cache[127][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27385_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01197_),
    .RESET_B(net322),
    .Q(\line_cache[127][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27386_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01198_),
    .RESET_B(net322),
    .Q(\line_cache[127][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27387_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01199_),
    .RESET_B(net322),
    .Q(\line_cache[127][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27388_ (.CLK(clknet_leaf_150_clk_i),
    .D(_01200_),
    .RESET_B(net312),
    .Q(\line_cache[127][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27389_ (.CLK(clknet_leaf_153_clk_i),
    .D(_01201_),
    .RESET_B(net322),
    .Q(\line_cache[127][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27390_ (.CLK(clknet_leaf_170_clk_i),
    .D(_01202_),
    .RESET_B(net323),
    .Q(\line_cache[127][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27391_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01203_),
    .RESET_B(net237),
    .Q(\line_cache[128][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27392_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01204_),
    .RESET_B(net316),
    .Q(\line_cache[128][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27393_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01205_),
    .RESET_B(net236),
    .Q(\line_cache[128][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27394_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01206_),
    .RESET_B(net236),
    .Q(\line_cache[128][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27395_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01207_),
    .RESET_B(net237),
    .Q(\line_cache[128][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27396_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01208_),
    .RESET_B(net236),
    .Q(\line_cache[128][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27397_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01209_),
    .RESET_B(net236),
    .Q(\line_cache[128][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27398_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01210_),
    .RESET_B(net237),
    .Q(\line_cache[128][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27399_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01211_),
    .RESET_B(net237),
    .Q(\line_cache[129][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27400_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01212_),
    .RESET_B(net316),
    .Q(\line_cache[129][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27401_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01213_),
    .RESET_B(net236),
    .Q(\line_cache[129][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27402_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01214_),
    .RESET_B(net316),
    .Q(\line_cache[129][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27403_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01215_),
    .RESET_B(net316),
    .Q(\line_cache[129][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27404_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01216_),
    .RESET_B(net316),
    .Q(\line_cache[129][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27405_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01217_),
    .RESET_B(net236),
    .Q(\line_cache[129][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27406_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01218_),
    .RESET_B(net236),
    .Q(\line_cache[129][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27407_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01219_),
    .RESET_B(net316),
    .Q(\line_cache[130][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27408_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01220_),
    .RESET_B(net316),
    .Q(\line_cache[130][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27409_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01221_),
    .RESET_B(net316),
    .Q(\line_cache[130][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27410_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01222_),
    .RESET_B(net316),
    .Q(\line_cache[130][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27411_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01223_),
    .RESET_B(net318),
    .Q(\line_cache[130][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27412_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01224_),
    .RESET_B(net316),
    .Q(\line_cache[130][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27413_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01225_),
    .RESET_B(net316),
    .Q(\line_cache[130][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27414_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01226_),
    .RESET_B(net318),
    .Q(\line_cache[130][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27415_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01227_),
    .RESET_B(net318),
    .Q(\line_cache[131][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27416_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01228_),
    .RESET_B(net317),
    .Q(\line_cache[131][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27417_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01229_),
    .RESET_B(net316),
    .Q(\line_cache[131][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27418_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01230_),
    .RESET_B(net316),
    .Q(\line_cache[131][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27419_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01231_),
    .RESET_B(net318),
    .Q(\line_cache[131][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27420_ (.CLK(clknet_leaf_157_clk_i),
    .D(_01232_),
    .RESET_B(net316),
    .Q(\line_cache[131][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27421_ (.CLK(clknet_leaf_156_clk_i),
    .D(_01233_),
    .RESET_B(net316),
    .Q(\line_cache[131][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27422_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01234_),
    .RESET_B(net318),
    .Q(\line_cache[131][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27423_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01235_),
    .RESET_B(net318),
    .Q(\line_cache[132][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27424_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01236_),
    .RESET_B(net320),
    .Q(\line_cache[132][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27425_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01237_),
    .RESET_B(net320),
    .Q(\line_cache[132][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27426_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01238_),
    .RESET_B(net320),
    .Q(\line_cache[132][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27427_ (.CLK(clknet_leaf_163_clk_i),
    .D(_01239_),
    .RESET_B(net320),
    .Q(\line_cache[132][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27428_ (.CLK(clknet_leaf_163_clk_i),
    .D(_01240_),
    .RESET_B(net320),
    .Q(\line_cache[132][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27429_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01241_),
    .RESET_B(net320),
    .Q(\line_cache[132][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27430_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01242_),
    .RESET_B(net320),
    .Q(\line_cache[132][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27431_ (.CLK(clknet_leaf_154_clk_i),
    .D(_01243_),
    .RESET_B(net323),
    .Q(\line_cache[133][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27432_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01244_),
    .RESET_B(net326),
    .Q(\line_cache[133][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27433_ (.CLK(clknet_leaf_165_clk_i),
    .D(_01245_),
    .RESET_B(net326),
    .Q(\line_cache[133][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27434_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01246_),
    .RESET_B(net326),
    .Q(\line_cache[133][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27435_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01247_),
    .RESET_B(net321),
    .Q(\line_cache[133][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27436_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01248_),
    .RESET_B(net326),
    .Q(\line_cache[133][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27437_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01249_),
    .RESET_B(net326),
    .Q(\line_cache[133][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27438_ (.CLK(clknet_leaf_165_clk_i),
    .D(_01250_),
    .RESET_B(net320),
    .Q(\line_cache[133][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27439_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01251_),
    .RESET_B(net320),
    .Q(\line_cache[134][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27440_ (.CLK(clknet_leaf_165_clk_i),
    .D(_01252_),
    .RESET_B(net326),
    .Q(\line_cache[134][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27441_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01253_),
    .RESET_B(net326),
    .Q(\line_cache[134][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27442_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01254_),
    .RESET_B(net320),
    .Q(\line_cache[134][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27443_ (.CLK(clknet_leaf_163_clk_i),
    .D(_01255_),
    .RESET_B(net321),
    .Q(\line_cache[134][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27444_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01256_),
    .RESET_B(net326),
    .Q(\line_cache[134][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27445_ (.CLK(clknet_leaf_170_clk_i),
    .D(_01257_),
    .RESET_B(net323),
    .Q(\line_cache[134][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27446_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01258_),
    .RESET_B(net327),
    .Q(\line_cache[134][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27447_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01259_),
    .RESET_B(net320),
    .Q(\line_cache[135][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27448_ (.CLK(clknet_leaf_165_clk_i),
    .D(_01260_),
    .RESET_B(net326),
    .Q(\line_cache[135][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27449_ (.CLK(clknet_leaf_169_clk_i),
    .D(_01261_),
    .RESET_B(net326),
    .Q(\line_cache[135][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27450_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01262_),
    .RESET_B(net320),
    .Q(\line_cache[135][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27451_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01263_),
    .RESET_B(net327),
    .Q(\line_cache[135][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27452_ (.CLK(clknet_leaf_166_clk_i),
    .D(_01264_),
    .RESET_B(net327),
    .Q(\line_cache[135][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27453_ (.CLK(clknet_leaf_170_clk_i),
    .D(_01265_),
    .RESET_B(net323),
    .Q(\line_cache[135][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27454_ (.CLK(clknet_leaf_165_clk_i),
    .D(_01266_),
    .RESET_B(net326),
    .Q(\line_cache[135][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27455_ (.CLK(clknet_leaf_158_clk_i),
    .D(_01267_),
    .RESET_B(net318),
    .Q(\line_cache[136][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27456_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01268_),
    .RESET_B(net319),
    .Q(\line_cache[136][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27457_ (.CLK(clknet_leaf_163_clk_i),
    .D(_01269_),
    .RESET_B(net321),
    .Q(\line_cache[136][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27458_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01270_),
    .RESET_B(net320),
    .Q(\line_cache[136][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27459_ (.CLK(clknet_leaf_163_clk_i),
    .D(_01271_),
    .RESET_B(net321),
    .Q(\line_cache[136][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27460_ (.CLK(clknet_leaf_163_clk_i),
    .D(_01272_),
    .RESET_B(net321),
    .Q(\line_cache[136][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27461_ (.CLK(clknet_leaf_159_clk_i),
    .D(_01273_),
    .RESET_B(net320),
    .Q(\line_cache[136][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27462_ (.CLK(clknet_leaf_164_clk_i),
    .D(_01274_),
    .RESET_B(net320),
    .Q(\line_cache[136][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27463_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01275_),
    .RESET_B(net319),
    .Q(\line_cache[137][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27464_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01276_),
    .RESET_B(net319),
    .Q(\line_cache[137][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27465_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01277_),
    .RESET_B(net319),
    .Q(\line_cache[137][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27466_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01278_),
    .RESET_B(net320),
    .Q(\line_cache[137][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27467_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01279_),
    .RESET_B(net321),
    .Q(\line_cache[137][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27468_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01280_),
    .RESET_B(net321),
    .Q(\line_cache[137][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27469_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01281_),
    .RESET_B(net319),
    .Q(\line_cache[137][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27470_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01282_),
    .RESET_B(net319),
    .Q(\line_cache[137][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27471_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01283_),
    .RESET_B(net319),
    .Q(\line_cache[138][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27472_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01284_),
    .RESET_B(net319),
    .Q(\line_cache[138][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27473_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01285_),
    .RESET_B(net319),
    .Q(\line_cache[138][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27474_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01286_),
    .RESET_B(net319),
    .Q(\line_cache[138][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27475_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01287_),
    .RESET_B(net319),
    .Q(\line_cache[138][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27476_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01288_),
    .RESET_B(net321),
    .Q(\line_cache[138][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27477_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01289_),
    .RESET_B(net319),
    .Q(\line_cache[138][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27478_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01290_),
    .RESET_B(net319),
    .Q(\line_cache[138][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27479_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01291_),
    .RESET_B(net318),
    .Q(\line_cache[139][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27480_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01292_),
    .RESET_B(net321),
    .Q(\line_cache[139][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27481_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01293_),
    .RESET_B(net321),
    .Q(\line_cache[139][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27482_ (.CLK(clknet_leaf_160_clk_i),
    .D(_01294_),
    .RESET_B(net319),
    .Q(\line_cache[139][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27483_ (.CLK(clknet_leaf_162_clk_i),
    .D(_01295_),
    .RESET_B(net321),
    .Q(\line_cache[139][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27484_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01296_),
    .RESET_B(net321),
    .Q(\line_cache[139][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27485_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01297_),
    .RESET_B(net319),
    .Q(\line_cache[139][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27486_ (.CLK(clknet_leaf_161_clk_i),
    .D(_01298_),
    .RESET_B(net319),
    .Q(\line_cache[139][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27487_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01299_),
    .RESET_B(net240),
    .Q(\line_cache[140][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27488_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01300_),
    .RESET_B(net240),
    .Q(\line_cache[140][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27489_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01301_),
    .RESET_B(net238),
    .Q(\line_cache[140][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27490_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01302_),
    .RESET_B(net240),
    .Q(\line_cache[140][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27491_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01303_),
    .RESET_B(net238),
    .Q(\line_cache[140][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27492_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01304_),
    .RESET_B(net238),
    .Q(\line_cache[140][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27493_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01305_),
    .RESET_B(net237),
    .Q(\line_cache[140][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27494_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01306_),
    .RESET_B(net237),
    .Q(\line_cache[140][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27495_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01307_),
    .RESET_B(net240),
    .Q(\line_cache[141][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27496_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01308_),
    .RESET_B(net240),
    .Q(\line_cache[141][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27497_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01309_),
    .RESET_B(net238),
    .Q(\line_cache[141][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27498_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01310_),
    .RESET_B(net240),
    .Q(\line_cache[141][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27499_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01311_),
    .RESET_B(net238),
    .Q(\line_cache[141][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27500_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01312_),
    .RESET_B(net239),
    .Q(\line_cache[141][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27501_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01313_),
    .RESET_B(net237),
    .Q(\line_cache[141][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27502_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01314_),
    .RESET_B(net237),
    .Q(\line_cache[141][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27503_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01315_),
    .RESET_B(net321),
    .Q(\line_cache[142][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27504_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01316_),
    .RESET_B(net241),
    .Q(\line_cache[142][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27505_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01317_),
    .RESET_B(net241),
    .Q(\line_cache[142][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27506_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01318_),
    .RESET_B(net240),
    .Q(\line_cache[142][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27507_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01319_),
    .RESET_B(net241),
    .Q(\line_cache[142][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27508_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01320_),
    .RESET_B(net241),
    .Q(\line_cache[142][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27509_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01321_),
    .RESET_B(net240),
    .Q(\line_cache[142][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27510_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01322_),
    .RESET_B(net240),
    .Q(\line_cache[142][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27511_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01323_),
    .RESET_B(net241),
    .Q(\line_cache[143][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27512_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01324_),
    .RESET_B(net321),
    .Q(\line_cache[143][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27513_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01325_),
    .RESET_B(net240),
    .Q(\line_cache[143][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27514_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01326_),
    .RESET_B(net240),
    .Q(\line_cache[143][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27515_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01327_),
    .RESET_B(net241),
    .Q(\line_cache[143][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27516_ (.CLK(clknet_leaf_116_clk_i),
    .D(_01328_),
    .RESET_B(net241),
    .Q(\line_cache[143][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27517_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01329_),
    .RESET_B(net240),
    .Q(\line_cache[143][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27518_ (.CLK(clknet_leaf_117_clk_i),
    .D(_01330_),
    .RESET_B(net240),
    .Q(\line_cache[143][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27519_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01331_),
    .RESET_B(net229),
    .Q(\line_cache[144][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27520_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01332_),
    .RESET_B(net236),
    .Q(\line_cache[144][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27521_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01333_),
    .RESET_B(net229),
    .Q(\line_cache[144][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27522_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01334_),
    .RESET_B(net235),
    .Q(\line_cache[144][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27523_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01335_),
    .RESET_B(net235),
    .Q(\line_cache[144][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27524_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01336_),
    .RESET_B(net236),
    .Q(\line_cache[144][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27525_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01337_),
    .RESET_B(net235),
    .Q(\line_cache[144][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27526_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01338_),
    .RESET_B(net235),
    .Q(\line_cache[144][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27527_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01339_),
    .RESET_B(net229),
    .Q(\line_cache[145][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27528_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01340_),
    .RESET_B(net236),
    .Q(\line_cache[145][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27529_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01341_),
    .RESET_B(net229),
    .Q(\line_cache[145][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27530_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01342_),
    .RESET_B(net235),
    .Q(\line_cache[145][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27531_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01343_),
    .RESET_B(net229),
    .Q(\line_cache[145][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27532_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01344_),
    .RESET_B(net236),
    .Q(\line_cache[145][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27533_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01345_),
    .RESET_B(net235),
    .Q(\line_cache[145][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27534_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01346_),
    .RESET_B(net235),
    .Q(\line_cache[145][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27535_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01347_),
    .RESET_B(net219),
    .Q(\line_cache[146][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27536_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01348_),
    .RESET_B(net236),
    .Q(\line_cache[146][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27537_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01349_),
    .RESET_B(net219),
    .Q(\line_cache[146][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27538_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01350_),
    .RESET_B(net235),
    .Q(\line_cache[146][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27539_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01351_),
    .RESET_B(net229),
    .Q(\line_cache[146][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27540_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01352_),
    .RESET_B(net235),
    .Q(\line_cache[146][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27541_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01353_),
    .RESET_B(net225),
    .Q(\line_cache[146][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27542_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01354_),
    .RESET_B(net225),
    .Q(\line_cache[146][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27543_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01355_),
    .RESET_B(net220),
    .Q(\line_cache[147][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27544_ (.CLK(clknet_leaf_121_clk_i),
    .D(_01356_),
    .RESET_B(net236),
    .Q(\line_cache[147][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27545_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01357_),
    .RESET_B(net225),
    .Q(\line_cache[147][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27546_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01358_),
    .RESET_B(net235),
    .Q(\line_cache[147][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27547_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01359_),
    .RESET_B(net235),
    .Q(\line_cache[147][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27548_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01360_),
    .RESET_B(net236),
    .Q(\line_cache[147][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27549_ (.CLK(clknet_leaf_133_clk_i),
    .D(_01361_),
    .RESET_B(net225),
    .Q(\line_cache[147][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27550_ (.CLK(clknet_leaf_122_clk_i),
    .D(_01362_),
    .RESET_B(net225),
    .Q(\line_cache[147][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27551_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01363_),
    .RESET_B(net240),
    .Q(\line_cache[148][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27552_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01364_),
    .RESET_B(net237),
    .Q(\line_cache[148][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27553_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01365_),
    .RESET_B(net238),
    .Q(\line_cache[148][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27554_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01366_),
    .RESET_B(net235),
    .Q(\line_cache[148][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27555_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01367_),
    .RESET_B(net235),
    .Q(\line_cache[148][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27556_ (.CLK(clknet_leaf_120_clk_i),
    .D(_01368_),
    .RESET_B(net237),
    .Q(\line_cache[148][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27557_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01369_),
    .RESET_B(net238),
    .Q(\line_cache[148][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27558_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01370_),
    .RESET_B(net235),
    .Q(\line_cache[148][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27559_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01371_),
    .RESET_B(net240),
    .Q(\line_cache[149][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27560_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01372_),
    .RESET_B(net237),
    .Q(\line_cache[149][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27561_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01373_),
    .RESET_B(net238),
    .Q(\line_cache[149][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27562_ (.CLK(clknet_leaf_123_clk_i),
    .D(_01374_),
    .RESET_B(net235),
    .Q(\line_cache[149][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27563_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01375_),
    .RESET_B(net235),
    .Q(\line_cache[149][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27564_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01376_),
    .RESET_B(net237),
    .Q(\line_cache[149][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27565_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01377_),
    .RESET_B(net238),
    .Q(\line_cache[149][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27566_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01378_),
    .RESET_B(net242),
    .Q(\line_cache[149][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27567_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01379_),
    .RESET_B(net238),
    .Q(\line_cache[150][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27568_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01380_),
    .RESET_B(net238),
    .Q(\line_cache[150][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27569_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01381_),
    .RESET_B(net239),
    .Q(\line_cache[150][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27570_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01382_),
    .RESET_B(net238),
    .Q(\line_cache[150][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27571_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01383_),
    .RESET_B(net242),
    .Q(\line_cache[150][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27572_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01384_),
    .RESET_B(net237),
    .Q(\line_cache[150][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27573_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01385_),
    .RESET_B(net239),
    .Q(\line_cache[150][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27574_ (.CLK(clknet_leaf_119_clk_i),
    .D(_01386_),
    .RESET_B(net242),
    .Q(\line_cache[150][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27575_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01387_),
    .RESET_B(net239),
    .Q(\line_cache[151][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27576_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01388_),
    .RESET_B(net238),
    .Q(\line_cache[151][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27577_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01389_),
    .RESET_B(net239),
    .Q(\line_cache[151][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27578_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01390_),
    .RESET_B(net238),
    .Q(\line_cache[151][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27579_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01391_),
    .RESET_B(net238),
    .Q(\line_cache[151][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27580_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01392_),
    .RESET_B(net240),
    .Q(\line_cache[151][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27581_ (.CLK(clknet_leaf_114_clk_i),
    .D(_01393_),
    .RESET_B(net239),
    .Q(\line_cache[151][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27582_ (.CLK(clknet_leaf_118_clk_i),
    .D(_01394_),
    .RESET_B(net238),
    .Q(\line_cache[151][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27583_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01395_),
    .RESET_B(net233),
    .Q(\line_cache[152][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27584_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01396_),
    .RESET_B(net233),
    .Q(\line_cache[152][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27585_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01397_),
    .RESET_B(net233),
    .Q(\line_cache[152][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27586_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01398_),
    .RESET_B(net231),
    .Q(\line_cache[152][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27587_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01399_),
    .RESET_B(net231),
    .Q(\line_cache[152][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27588_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01400_),
    .RESET_B(net233),
    .Q(\line_cache[152][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27589_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01401_),
    .RESET_B(net233),
    .Q(\line_cache[152][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27590_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01402_),
    .RESET_B(net233),
    .Q(\line_cache[152][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27591_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01403_),
    .RESET_B(net239),
    .Q(\line_cache[153][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27592_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01404_),
    .RESET_B(net239),
    .Q(\line_cache[153][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27593_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01405_),
    .RESET_B(net234),
    .Q(\line_cache[153][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27594_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01406_),
    .RESET_B(net231),
    .Q(\line_cache[153][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27595_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01407_),
    .RESET_B(net231),
    .Q(\line_cache[153][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27596_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01408_),
    .RESET_B(net234),
    .Q(\line_cache[153][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27597_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01409_),
    .RESET_B(net233),
    .Q(\line_cache[153][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27598_ (.CLK(clknet_leaf_113_clk_i),
    .D(_01410_),
    .RESET_B(net233),
    .Q(\line_cache[153][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27599_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01411_),
    .RESET_B(net239),
    .Q(\line_cache[154][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27600_ (.CLK(clknet_leaf_115_clk_i),
    .D(_01412_),
    .RESET_B(net239),
    .Q(\line_cache[154][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27601_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01413_),
    .RESET_B(net231),
    .Q(\line_cache[154][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27602_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01414_),
    .RESET_B(net234),
    .Q(\line_cache[154][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27603_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01415_),
    .RESET_B(net234),
    .Q(\line_cache[154][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27604_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01416_),
    .RESET_B(net234),
    .Q(\line_cache[154][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27605_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01417_),
    .RESET_B(net234),
    .Q(\line_cache[154][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27606_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01418_),
    .RESET_B(net233),
    .Q(\line_cache[154][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27607_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01419_),
    .RESET_B(net234),
    .Q(\line_cache[155][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27608_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01420_),
    .RESET_B(net234),
    .Q(\line_cache[155][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27609_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01421_),
    .RESET_B(net234),
    .Q(\line_cache[155][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27610_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01422_),
    .RESET_B(net231),
    .Q(\line_cache[155][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27611_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01423_),
    .RESET_B(net232),
    .Q(\line_cache[155][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27612_ (.CLK(clknet_leaf_111_clk_i),
    .D(_01424_),
    .RESET_B(net234),
    .Q(\line_cache[155][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27613_ (.CLK(clknet_leaf_112_clk_i),
    .D(_01425_),
    .RESET_B(net233),
    .Q(\line_cache[155][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27614_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01426_),
    .RESET_B(net233),
    .Q(\line_cache[155][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27615_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01427_),
    .RESET_B(net233),
    .Q(\line_cache[156][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27616_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01428_),
    .RESET_B(net233),
    .Q(\line_cache[156][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27617_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01429_),
    .RESET_B(net231),
    .Q(\line_cache[156][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27618_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01430_),
    .RESET_B(net228),
    .Q(\line_cache[156][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27619_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01431_),
    .RESET_B(net228),
    .Q(\line_cache[156][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27620_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01432_),
    .RESET_B(net231),
    .Q(\line_cache[156][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27621_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01433_),
    .RESET_B(net233),
    .Q(\line_cache[156][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27622_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01434_),
    .RESET_B(net233),
    .Q(\line_cache[156][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27623_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01435_),
    .RESET_B(net233),
    .Q(\line_cache[157][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27624_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01436_),
    .RESET_B(net229),
    .Q(\line_cache[157][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27625_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01437_),
    .RESET_B(net228),
    .Q(\line_cache[157][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27626_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01438_),
    .RESET_B(net228),
    .Q(\line_cache[157][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27627_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01439_),
    .RESET_B(net228),
    .Q(\line_cache[157][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27628_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01440_),
    .RESET_B(net228),
    .Q(\line_cache[157][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27629_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01441_),
    .RESET_B(net231),
    .Q(\line_cache[157][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27630_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01442_),
    .RESET_B(net229),
    .Q(\line_cache[157][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27631_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01443_),
    .RESET_B(net229),
    .Q(\line_cache[158][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27632_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01444_),
    .RESET_B(net229),
    .Q(\line_cache[158][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27633_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01445_),
    .RESET_B(net230),
    .Q(\line_cache[158][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27634_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01446_),
    .RESET_B(net228),
    .Q(\line_cache[158][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27635_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01447_),
    .RESET_B(net230),
    .Q(\line_cache[158][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27636_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01448_),
    .RESET_B(net229),
    .Q(\line_cache[158][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27637_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01449_),
    .RESET_B(net230),
    .Q(\line_cache[158][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27638_ (.CLK(clknet_leaf_125_clk_i),
    .D(_01450_),
    .RESET_B(net229),
    .Q(\line_cache[158][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27639_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01451_),
    .RESET_B(net230),
    .Q(\line_cache[159][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27640_ (.CLK(clknet_leaf_124_clk_i),
    .D(_01452_),
    .RESET_B(net230),
    .Q(\line_cache[159][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27641_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01453_),
    .RESET_B(net230),
    .Q(\line_cache[159][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27642_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01454_),
    .RESET_B(net228),
    .Q(\line_cache[159][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27643_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01455_),
    .RESET_B(net209),
    .Q(\line_cache[159][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27644_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01456_),
    .RESET_B(net230),
    .Q(\line_cache[159][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27645_ (.CLK(clknet_leaf_105_clk_i),
    .D(_01457_),
    .RESET_B(net230),
    .Q(\line_cache[159][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27646_ (.CLK(clknet_leaf_106_clk_i),
    .D(_01458_),
    .RESET_B(net230),
    .Q(\line_cache[159][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27647_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01459_),
    .RESET_B(net207),
    .Q(\line_cache[160][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27648_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01460_),
    .RESET_B(net207),
    .Q(\line_cache[160][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27649_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01461_),
    .RESET_B(net202),
    .Q(\line_cache[160][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27650_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01462_),
    .RESET_B(net207),
    .Q(\line_cache[160][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27651_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01463_),
    .RESET_B(net203),
    .Q(\line_cache[160][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27652_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01464_),
    .RESET_B(net207),
    .Q(\line_cache[160][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27653_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01465_),
    .RESET_B(net207),
    .Q(\line_cache[160][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27654_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01466_),
    .RESET_B(net204),
    .Q(\line_cache[160][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27655_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01467_),
    .RESET_B(net207),
    .Q(\line_cache[161][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27656_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01468_),
    .RESET_B(net206),
    .Q(\line_cache[161][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27657_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01469_),
    .RESET_B(net203),
    .Q(\line_cache[161][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27658_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01470_),
    .RESET_B(net207),
    .Q(\line_cache[161][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27659_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01471_),
    .RESET_B(net203),
    .Q(\line_cache[161][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27660_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01472_),
    .RESET_B(net203),
    .Q(\line_cache[161][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27661_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01473_),
    .RESET_B(net207),
    .Q(\line_cache[161][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27662_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01474_),
    .RESET_B(net204),
    .Q(\line_cache[161][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27663_ (.CLK(clknet_leaf_92_clk_i),
    .D(_01475_),
    .RESET_B(net207),
    .Q(\line_cache[162][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27664_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01476_),
    .RESET_B(net204),
    .Q(\line_cache[162][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27665_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01477_),
    .RESET_B(net203),
    .Q(\line_cache[162][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27666_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01478_),
    .RESET_B(net204),
    .Q(\line_cache[162][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27667_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01479_),
    .RESET_B(net203),
    .Q(\line_cache[162][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27668_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01480_),
    .RESET_B(net203),
    .Q(\line_cache[162][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27669_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01481_),
    .RESET_B(net204),
    .Q(\line_cache[162][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27670_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01482_),
    .RESET_B(net208),
    .Q(\line_cache[162][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27671_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01483_),
    .RESET_B(net207),
    .Q(\line_cache[163][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27672_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01484_),
    .RESET_B(net204),
    .Q(\line_cache[163][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27673_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01485_),
    .RESET_B(net203),
    .Q(\line_cache[163][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27674_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01486_),
    .RESET_B(net204),
    .Q(\line_cache[163][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27675_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01487_),
    .RESET_B(net203),
    .Q(\line_cache[163][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27676_ (.CLK(clknet_leaf_88_clk_i),
    .D(_01488_),
    .RESET_B(net203),
    .Q(\line_cache[163][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27677_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01489_),
    .RESET_B(net208),
    .Q(\line_cache[163][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27678_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01490_),
    .RESET_B(net208),
    .Q(\line_cache[163][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27679_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01491_),
    .RESET_B(net206),
    .Q(\line_cache[164][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27680_ (.CLK(clknet_leaf_91_clk_i),
    .D(_01492_),
    .RESET_B(net207),
    .Q(\line_cache[164][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27681_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01493_),
    .RESET_B(net206),
    .Q(\line_cache[164][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27682_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01494_),
    .RESET_B(net204),
    .Q(\line_cache[164][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27683_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01495_),
    .RESET_B(net206),
    .Q(\line_cache[164][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27684_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01496_),
    .RESET_B(net206),
    .Q(\line_cache[164][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27685_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01497_),
    .RESET_B(net206),
    .Q(\line_cache[164][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27686_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01498_),
    .RESET_B(net204),
    .Q(\line_cache[164][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27687_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01499_),
    .RESET_B(net206),
    .Q(\line_cache[165][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27688_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01500_),
    .RESET_B(net206),
    .Q(\line_cache[165][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27689_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01501_),
    .RESET_B(net206),
    .Q(\line_cache[165][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27690_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01502_),
    .RESET_B(net205),
    .Q(\line_cache[165][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27691_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01503_),
    .RESET_B(net206),
    .Q(\line_cache[165][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27692_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01504_),
    .RESET_B(net205),
    .Q(\line_cache[165][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27693_ (.CLK(clknet_leaf_90_clk_i),
    .D(_01505_),
    .RESET_B(net206),
    .Q(\line_cache[165][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27694_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01506_),
    .RESET_B(net208),
    .Q(\line_cache[165][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27695_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01507_),
    .RESET_B(net206),
    .Q(\line_cache[166][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27696_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01508_),
    .RESET_B(net211),
    .Q(\line_cache[166][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27697_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01509_),
    .RESET_B(net211),
    .Q(\line_cache[166][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27698_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01510_),
    .RESET_B(net208),
    .Q(\line_cache[166][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27699_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01511_),
    .RESET_B(net211),
    .Q(\line_cache[166][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27700_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01512_),
    .RESET_B(net208),
    .Q(\line_cache[166][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27701_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01513_),
    .RESET_B(net211),
    .Q(\line_cache[166][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27702_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01514_),
    .RESET_B(net210),
    .Q(\line_cache[166][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27703_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01515_),
    .RESET_B(net211),
    .Q(\line_cache[167][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27704_ (.CLK(clknet_leaf_94_clk_i),
    .D(_01516_),
    .RESET_B(net206),
    .Q(\line_cache[167][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27705_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01517_),
    .RESET_B(net211),
    .Q(\line_cache[167][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27706_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01518_),
    .RESET_B(net210),
    .Q(\line_cache[167][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27707_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01519_),
    .RESET_B(net212),
    .Q(\line_cache[167][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27708_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01520_),
    .RESET_B(net209),
    .Q(\line_cache[167][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27709_ (.CLK(clknet_leaf_95_clk_i),
    .D(_01521_),
    .RESET_B(net211),
    .Q(\line_cache[167][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27710_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01522_),
    .RESET_B(net212),
    .Q(\line_cache[167][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27711_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01523_),
    .RESET_B(net212),
    .Q(\line_cache[168][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27712_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01524_),
    .RESET_B(net232),
    .Q(\line_cache[168][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27713_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01525_),
    .RESET_B(net232),
    .Q(\line_cache[168][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27714_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01526_),
    .RESET_B(net231),
    .Q(\line_cache[168][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27715_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01527_),
    .RESET_B(net212),
    .Q(\line_cache[168][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27716_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01528_),
    .RESET_B(net209),
    .Q(\line_cache[168][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27717_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01529_),
    .RESET_B(net209),
    .Q(\line_cache[168][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27718_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01530_),
    .RESET_B(net230),
    .Q(\line_cache[168][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27719_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01531_),
    .RESET_B(net212),
    .Q(\line_cache[169][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27720_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01532_),
    .RESET_B(net232),
    .Q(\line_cache[169][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27721_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01533_),
    .RESET_B(net232),
    .Q(\line_cache[169][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27722_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01534_),
    .RESET_B(net231),
    .Q(\line_cache[169][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27723_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01535_),
    .RESET_B(net212),
    .Q(\line_cache[169][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27724_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01536_),
    .RESET_B(net212),
    .Q(\line_cache[169][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27725_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01537_),
    .RESET_B(net212),
    .Q(\line_cache[169][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27726_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01538_),
    .RESET_B(net231),
    .Q(\line_cache[169][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27727_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01539_),
    .RESET_B(net212),
    .Q(\line_cache[170][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27728_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01540_),
    .RESET_B(net232),
    .Q(\line_cache[170][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27729_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01541_),
    .RESET_B(net232),
    .Q(\line_cache[170][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27730_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01542_),
    .RESET_B(net231),
    .Q(\line_cache[170][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27731_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01543_),
    .RESET_B(net212),
    .Q(\line_cache[170][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27732_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01544_),
    .RESET_B(net212),
    .Q(\line_cache[170][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27733_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01545_),
    .RESET_B(net212),
    .Q(\line_cache[170][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27734_ (.CLK(clknet_leaf_107_clk_i),
    .D(_01546_),
    .RESET_B(net231),
    .Q(\line_cache[170][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27735_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01547_),
    .RESET_B(net212),
    .Q(\line_cache[171][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27736_ (.CLK(clknet_leaf_109_clk_i),
    .D(_01548_),
    .RESET_B(net232),
    .Q(\line_cache[171][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27737_ (.CLK(clknet_leaf_110_clk_i),
    .D(_01549_),
    .RESET_B(net232),
    .Q(\line_cache[171][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27738_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01550_),
    .RESET_B(net231),
    .Q(\line_cache[171][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27739_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01551_),
    .RESET_B(net213),
    .Q(\line_cache[171][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27740_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01552_),
    .RESET_B(net212),
    .Q(\line_cache[171][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27741_ (.CLK(clknet_leaf_99_clk_i),
    .D(_01553_),
    .RESET_B(net212),
    .Q(\line_cache[171][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27742_ (.CLK(clknet_leaf_108_clk_i),
    .D(_01554_),
    .RESET_B(net231),
    .Q(\line_cache[171][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27743_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01555_),
    .RESET_B(net206),
    .Q(\line_cache[172][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27744_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01556_),
    .RESET_B(net211),
    .Q(\line_cache[172][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27745_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01557_),
    .RESET_B(net206),
    .Q(\line_cache[172][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27746_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01558_),
    .RESET_B(net206),
    .Q(\line_cache[172][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27747_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01559_),
    .RESET_B(net214),
    .Q(\line_cache[172][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27748_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01560_),
    .RESET_B(net211),
    .Q(\line_cache[172][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27749_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01561_),
    .RESET_B(net214),
    .Q(\line_cache[172][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27750_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01562_),
    .RESET_B(net214),
    .Q(\line_cache[172][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27751_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01563_),
    .RESET_B(net207),
    .Q(\line_cache[173][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27752_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01564_),
    .RESET_B(net211),
    .Q(\line_cache[173][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27753_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01565_),
    .RESET_B(net207),
    .Q(\line_cache[173][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27754_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01566_),
    .RESET_B(net212),
    .Q(\line_cache[173][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27755_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01567_),
    .RESET_B(net207),
    .Q(\line_cache[173][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27756_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01568_),
    .RESET_B(net213),
    .Q(\line_cache[173][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27757_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01569_),
    .RESET_B(net207),
    .Q(\line_cache[173][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27758_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01570_),
    .RESET_B(net211),
    .Q(\line_cache[173][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27759_ (.CLK(clknet_leaf_93_clk_i),
    .D(_01571_),
    .RESET_B(net211),
    .Q(\line_cache[174][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27760_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01572_),
    .RESET_B(net211),
    .Q(\line_cache[174][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27761_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01573_),
    .RESET_B(net211),
    .Q(\line_cache[174][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27762_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01574_),
    .RESET_B(net213),
    .Q(\line_cache[174][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27763_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01575_),
    .RESET_B(net211),
    .Q(\line_cache[174][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27764_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01576_),
    .RESET_B(net213),
    .Q(\line_cache[174][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27765_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01577_),
    .RESET_B(net211),
    .Q(\line_cache[174][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27766_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01578_),
    .RESET_B(net213),
    .Q(\line_cache[174][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27767_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01579_),
    .RESET_B(net213),
    .Q(\line_cache[175][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27768_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01580_),
    .RESET_B(net213),
    .Q(\line_cache[175][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27769_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01581_),
    .RESET_B(net213),
    .Q(\line_cache[175][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27770_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01582_),
    .RESET_B(net213),
    .Q(\line_cache[175][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27771_ (.CLK(clknet_leaf_97_clk_i),
    .D(_01583_),
    .RESET_B(net213),
    .Q(\line_cache[175][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27772_ (.CLK(clknet_leaf_98_clk_i),
    .D(_01584_),
    .RESET_B(net213),
    .Q(\line_cache[175][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27773_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01585_),
    .RESET_B(net213),
    .Q(\line_cache[175][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27774_ (.CLK(clknet_leaf_96_clk_i),
    .D(_01586_),
    .RESET_B(net213),
    .Q(\line_cache[175][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27775_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01587_),
    .RESET_B(net203),
    .Q(\line_cache[176][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27776_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01588_),
    .RESET_B(net203),
    .Q(\line_cache[176][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27777_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01589_),
    .RESET_B(net202),
    .Q(\line_cache[176][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27778_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01590_),
    .RESET_B(net202),
    .Q(\line_cache[176][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27779_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01591_),
    .RESET_B(net202),
    .Q(\line_cache[176][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27780_ (.CLK(clknet_leaf_87_clk_i),
    .D(_01592_),
    .RESET_B(net202),
    .Q(\line_cache[176][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27781_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01593_),
    .RESET_B(net202),
    .Q(\line_cache[176][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27782_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01594_),
    .RESET_B(net202),
    .Q(\line_cache[176][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27783_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01595_),
    .RESET_B(net202),
    .Q(\line_cache[177][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27784_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01596_),
    .RESET_B(net202),
    .Q(\line_cache[177][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27785_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01597_),
    .RESET_B(net202),
    .Q(\line_cache[177][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27786_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01598_),
    .RESET_B(net202),
    .Q(\line_cache[177][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27787_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01599_),
    .RESET_B(net202),
    .Q(\line_cache[177][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27788_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01600_),
    .RESET_B(net202),
    .Q(\line_cache[177][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27789_ (.CLK(clknet_leaf_86_clk_i),
    .D(_01601_),
    .RESET_B(net202),
    .Q(\line_cache[177][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27790_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01602_),
    .RESET_B(net202),
    .Q(\line_cache[177][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27791_ (.CLK(clknet_leaf_89_clk_i),
    .D(_01603_),
    .RESET_B(net205),
    .Q(\line_cache[178][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27792_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01604_),
    .RESET_B(net204),
    .Q(\line_cache[178][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27793_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01605_),
    .RESET_B(net202),
    .Q(\line_cache[178][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27794_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01606_),
    .RESET_B(net204),
    .Q(\line_cache[178][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27795_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01607_),
    .RESET_B(net204),
    .Q(\line_cache[178][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27796_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01608_),
    .RESET_B(net210),
    .Q(\line_cache[178][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27797_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01609_),
    .RESET_B(net192),
    .Q(\line_cache[178][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27798_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01610_),
    .RESET_B(net208),
    .Q(\line_cache[178][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27799_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01611_),
    .RESET_B(net205),
    .Q(\line_cache[179][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27800_ (.CLK(clknet_leaf_84_clk_i),
    .D(_01612_),
    .RESET_B(net205),
    .Q(\line_cache[179][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27801_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01613_),
    .RESET_B(net204),
    .Q(\line_cache[179][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27802_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01614_),
    .RESET_B(net204),
    .Q(\line_cache[179][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27803_ (.CLK(clknet_leaf_85_clk_i),
    .D(_01615_),
    .RESET_B(net204),
    .Q(\line_cache[179][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27804_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01616_),
    .RESET_B(net208),
    .Q(\line_cache[179][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27805_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01617_),
    .RESET_B(net204),
    .Q(\line_cache[179][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27806_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01618_),
    .RESET_B(net208),
    .Q(\line_cache[179][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27807_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01619_),
    .RESET_B(net228),
    .Q(\line_cache[180][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27808_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01620_),
    .RESET_B(net228),
    .Q(\line_cache[180][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27809_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01621_),
    .RESET_B(net220),
    .Q(\line_cache[180][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27810_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01622_),
    .RESET_B(net228),
    .Q(\line_cache[180][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27811_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01623_),
    .RESET_B(net218),
    .Q(\line_cache[180][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27812_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01624_),
    .RESET_B(net220),
    .Q(\line_cache[180][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27813_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01625_),
    .RESET_B(net220),
    .Q(\line_cache[180][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27814_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01626_),
    .RESET_B(net228),
    .Q(\line_cache[180][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27815_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01627_),
    .RESET_B(net228),
    .Q(\line_cache[181][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27816_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01628_),
    .RESET_B(net228),
    .Q(\line_cache[181][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27817_ (.CLK(clknet_leaf_130_clk_i),
    .D(_01629_),
    .RESET_B(net220),
    .Q(\line_cache[181][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27818_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01630_),
    .RESET_B(net218),
    .Q(\line_cache[181][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27819_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01631_),
    .RESET_B(net218),
    .Q(\line_cache[181][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27820_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01632_),
    .RESET_B(net229),
    .Q(\line_cache[181][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27821_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01633_),
    .RESET_B(net218),
    .Q(\line_cache[181][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27822_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01634_),
    .RESET_B(net218),
    .Q(\line_cache[181][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27823_ (.CLK(clknet_leaf_104_clk_i),
    .D(_01635_),
    .RESET_B(net228),
    .Q(\line_cache[182][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27824_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01636_),
    .RESET_B(net209),
    .Q(\line_cache[182][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27825_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01637_),
    .RESET_B(net220),
    .Q(\line_cache[182][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27826_ (.CLK(clknet_leaf_81_clk_i),
    .D(_01638_),
    .RESET_B(net199),
    .Q(\line_cache[182][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27827_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01639_),
    .RESET_B(net218),
    .Q(\line_cache[182][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27828_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01640_),
    .RESET_B(net229),
    .Q(\line_cache[182][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27829_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01641_),
    .RESET_B(net221),
    .Q(\line_cache[182][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27830_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01642_),
    .RESET_B(net221),
    .Q(\line_cache[182][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27831_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01643_),
    .RESET_B(net229),
    .Q(\line_cache[183][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27832_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01644_),
    .RESET_B(net209),
    .Q(\line_cache[183][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27833_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01645_),
    .RESET_B(net220),
    .Q(\line_cache[183][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27834_ (.CLK(clknet_leaf_103_clk_i),
    .D(_01646_),
    .RESET_B(net209),
    .Q(\line_cache[183][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27835_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01647_),
    .RESET_B(net199),
    .Q(\line_cache[183][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27836_ (.CLK(clknet_leaf_126_clk_i),
    .D(_01648_),
    .RESET_B(net229),
    .Q(\line_cache[183][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27837_ (.CLK(clknet_leaf_128_clk_i),
    .D(_01649_),
    .RESET_B(net221),
    .Q(\line_cache[183][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27838_ (.CLK(clknet_leaf_127_clk_i),
    .D(_01650_),
    .RESET_B(net228),
    .Q(\line_cache[183][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27839_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01651_),
    .RESET_B(net190),
    .Q(\line_cache[184][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27840_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01652_),
    .RESET_B(net190),
    .Q(\line_cache[184][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27841_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01653_),
    .RESET_B(net190),
    .Q(\line_cache[184][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27842_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01654_),
    .RESET_B(net190),
    .Q(\line_cache[184][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27843_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01655_),
    .RESET_B(net190),
    .Q(\line_cache[184][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27844_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01656_),
    .RESET_B(net190),
    .Q(\line_cache[184][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27845_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01657_),
    .RESET_B(net190),
    .Q(\line_cache[184][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27846_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01658_),
    .RESET_B(net198),
    .Q(\line_cache[184][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27847_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01659_),
    .RESET_B(net191),
    .Q(\line_cache[185][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27848_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01660_),
    .RESET_B(net192),
    .Q(\line_cache[185][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27849_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01661_),
    .RESET_B(net191),
    .Q(\line_cache[185][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27850_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01662_),
    .RESET_B(net191),
    .Q(\line_cache[185][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27851_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01663_),
    .RESET_B(net191),
    .Q(\line_cache[185][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27852_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01664_),
    .RESET_B(net191),
    .Q(\line_cache[185][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27853_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01665_),
    .RESET_B(net192),
    .Q(\line_cache[185][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27854_ (.CLK(clknet_leaf_76_clk_i),
    .D(_01666_),
    .RESET_B(net192),
    .Q(\line_cache[185][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27855_ (.CLK(clknet_leaf_74_clk_i),
    .D(_01667_),
    .RESET_B(net191),
    .Q(\line_cache[186][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27856_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01668_),
    .RESET_B(net192),
    .Q(\line_cache[186][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27857_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01669_),
    .RESET_B(net190),
    .Q(\line_cache[186][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27858_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01670_),
    .RESET_B(net193),
    .Q(\line_cache[186][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27859_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01671_),
    .RESET_B(net191),
    .Q(\line_cache[186][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27860_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01672_),
    .RESET_B(net193),
    .Q(\line_cache[186][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27861_ (.CLK(clknet_leaf_76_clk_i),
    .D(_01673_),
    .RESET_B(net193),
    .Q(\line_cache[186][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27862_ (.CLK(clknet_leaf_76_clk_i),
    .D(_01674_),
    .RESET_B(net193),
    .Q(\line_cache[186][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27863_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01675_),
    .RESET_B(net191),
    .Q(\line_cache[187][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27864_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01676_),
    .RESET_B(net192),
    .Q(\line_cache[187][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27865_ (.CLK(clknet_leaf_73_clk_i),
    .D(_01677_),
    .RESET_B(net191),
    .Q(\line_cache[187][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27866_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01678_),
    .RESET_B(net193),
    .Q(\line_cache[187][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27867_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01679_),
    .RESET_B(net191),
    .Q(\line_cache[187][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27868_ (.CLK(clknet_leaf_75_clk_i),
    .D(_01680_),
    .RESET_B(net193),
    .Q(\line_cache[187][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27869_ (.CLK(clknet_leaf_76_clk_i),
    .D(_01681_),
    .RESET_B(net193),
    .Q(\line_cache[187][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27870_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01682_),
    .RESET_B(net198),
    .Q(\line_cache[187][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27871_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01683_),
    .RESET_B(net210),
    .Q(\line_cache[188][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27872_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01684_),
    .RESET_B(net209),
    .Q(\line_cache[188][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27873_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01685_),
    .RESET_B(net200),
    .Q(\line_cache[188][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27874_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01686_),
    .RESET_B(net208),
    .Q(\line_cache[188][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27875_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01687_),
    .RESET_B(net208),
    .Q(\line_cache[188][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27876_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01688_),
    .RESET_B(net209),
    .Q(\line_cache[188][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27877_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01689_),
    .RESET_B(net198),
    .Q(\line_cache[188][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27878_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01690_),
    .RESET_B(net208),
    .Q(\line_cache[188][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27879_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01691_),
    .RESET_B(net210),
    .Q(\line_cache[189][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27880_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01692_),
    .RESET_B(net210),
    .Q(\line_cache[189][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27881_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01693_),
    .RESET_B(net200),
    .Q(\line_cache[189][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27882_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01694_),
    .RESET_B(net208),
    .Q(\line_cache[189][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27883_ (.CLK(clknet_leaf_81_clk_i),
    .D(_01695_),
    .RESET_B(net209),
    .Q(\line_cache[189][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27884_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01696_),
    .RESET_B(net210),
    .Q(\line_cache[189][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27885_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01697_),
    .RESET_B(net198),
    .Q(\line_cache[189][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27886_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01698_),
    .RESET_B(net208),
    .Q(\line_cache[189][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27887_ (.CLK(clknet_leaf_83_clk_i),
    .D(_01699_),
    .RESET_B(net210),
    .Q(\line_cache[190][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27888_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01700_),
    .RESET_B(net210),
    .Q(\line_cache[190][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27889_ (.CLK(clknet_leaf_81_clk_i),
    .D(_01701_),
    .RESET_B(net209),
    .Q(\line_cache[190][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27890_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01702_),
    .RESET_B(net208),
    .Q(\line_cache[190][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27891_ (.CLK(clknet_leaf_81_clk_i),
    .D(_01703_),
    .RESET_B(net209),
    .Q(\line_cache[190][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27892_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01704_),
    .RESET_B(net210),
    .Q(\line_cache[190][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27893_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01705_),
    .RESET_B(net198),
    .Q(\line_cache[190][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27894_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01706_),
    .RESET_B(net209),
    .Q(\line_cache[190][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27895_ (.CLK(clknet_leaf_100_clk_i),
    .D(_01707_),
    .RESET_B(net210),
    .Q(\line_cache[191][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27896_ (.CLK(clknet_leaf_101_clk_i),
    .D(_01708_),
    .RESET_B(net210),
    .Q(\line_cache[191][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27897_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01709_),
    .RESET_B(net200),
    .Q(\line_cache[191][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27898_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01710_),
    .RESET_B(net209),
    .Q(\line_cache[191][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27899_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01711_),
    .RESET_B(net209),
    .Q(\line_cache[191][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27900_ (.CLK(clknet_leaf_102_clk_i),
    .D(_01712_),
    .RESET_B(net209),
    .Q(\line_cache[191][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27901_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01713_),
    .RESET_B(net198),
    .Q(\line_cache[191][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27902_ (.CLK(clknet_leaf_82_clk_i),
    .D(_01714_),
    .RESET_B(net208),
    .Q(\line_cache[191][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27903_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01715_),
    .RESET_B(net156),
    .Q(\line_cache[192][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27904_ (.CLK(clknet_leaf_31_clk_i),
    .D(_01716_),
    .RESET_B(net153),
    .Q(\line_cache[192][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27905_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01717_),
    .RESET_B(net156),
    .Q(\line_cache[192][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27906_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01718_),
    .RESET_B(net178),
    .Q(\line_cache[192][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27907_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01719_),
    .RESET_B(net175),
    .Q(\line_cache[192][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27908_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01720_),
    .RESET_B(net153),
    .Q(\line_cache[192][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27909_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01721_),
    .RESET_B(net156),
    .Q(\line_cache[192][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27910_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01722_),
    .RESET_B(net178),
    .Q(\line_cache[192][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27911_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01723_),
    .RESET_B(net156),
    .Q(\line_cache[193][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27912_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01724_),
    .RESET_B(net153),
    .Q(\line_cache[193][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27913_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01725_),
    .RESET_B(net156),
    .Q(\line_cache[193][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27914_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01726_),
    .RESET_B(net156),
    .Q(\line_cache[193][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27915_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01727_),
    .RESET_B(net153),
    .Q(\line_cache[193][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27916_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01728_),
    .RESET_B(net156),
    .Q(\line_cache[193][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27917_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01729_),
    .RESET_B(net156),
    .Q(\line_cache[193][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27918_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01730_),
    .RESET_B(net156),
    .Q(\line_cache[193][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27919_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01731_),
    .RESET_B(net156),
    .Q(\line_cache[194][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27920_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01732_),
    .RESET_B(net153),
    .Q(\line_cache[194][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27921_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01733_),
    .RESET_B(net156),
    .Q(\line_cache[194][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27922_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01734_),
    .RESET_B(net156),
    .Q(\line_cache[194][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27923_ (.CLK(clknet_leaf_28_clk_i),
    .D(_01735_),
    .RESET_B(net153),
    .Q(\line_cache[194][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27924_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01736_),
    .RESET_B(net156),
    .Q(\line_cache[194][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27925_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01737_),
    .RESET_B(net156),
    .Q(\line_cache[194][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27926_ (.CLK(clknet_leaf_26_clk_i),
    .D(_01738_),
    .RESET_B(net156),
    .Q(\line_cache[194][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27927_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01739_),
    .RESET_B(net155),
    .Q(\line_cache[195][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27928_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01740_),
    .RESET_B(net152),
    .Q(\line_cache[195][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27929_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01741_),
    .RESET_B(net155),
    .Q(\line_cache[195][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27930_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01742_),
    .RESET_B(net155),
    .Q(\line_cache[195][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27931_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01743_),
    .RESET_B(net152),
    .Q(\line_cache[195][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27932_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01744_),
    .RESET_B(net152),
    .Q(\line_cache[195][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27933_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01745_),
    .RESET_B(net155),
    .Q(\line_cache[195][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27934_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01746_),
    .RESET_B(net155),
    .Q(\line_cache[195][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27935_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01747_),
    .RESET_B(net155),
    .Q(\line_cache[196][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27936_ (.CLK(clknet_leaf_11_clk_i),
    .D(_01748_),
    .RESET_B(net152),
    .Q(\line_cache[196][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27937_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01749_),
    .RESET_B(net155),
    .Q(\line_cache[196][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27938_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01750_),
    .RESET_B(net155),
    .Q(\line_cache[196][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27939_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01751_),
    .RESET_B(net152),
    .Q(\line_cache[196][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27940_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01752_),
    .RESET_B(net152),
    .Q(\line_cache[196][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27941_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01753_),
    .RESET_B(net155),
    .Q(\line_cache[196][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27942_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01754_),
    .RESET_B(net155),
    .Q(\line_cache[196][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27943_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01755_),
    .RESET_B(net157),
    .Q(\line_cache[197][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27944_ (.CLK(clknet_leaf_11_clk_i),
    .D(_01756_),
    .RESET_B(net152),
    .Q(\line_cache[197][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27945_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01757_),
    .RESET_B(net157),
    .Q(\line_cache[197][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27946_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01758_),
    .RESET_B(net155),
    .Q(\line_cache[197][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27947_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01759_),
    .RESET_B(net150),
    .Q(\line_cache[197][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27948_ (.CLK(clknet_leaf_11_clk_i),
    .D(_01760_),
    .RESET_B(net152),
    .Q(\line_cache[197][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27949_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01761_),
    .RESET_B(net155),
    .Q(\line_cache[197][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27950_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01762_),
    .RESET_B(net155),
    .Q(\line_cache[197][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27951_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01763_),
    .RESET_B(net149),
    .Q(\line_cache[198][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27952_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01764_),
    .RESET_B(net149),
    .Q(\line_cache[198][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27953_ (.CLK(clknet_leaf_23_clk_i),
    .D(_01765_),
    .RESET_B(net157),
    .Q(\line_cache[198][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27954_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01766_),
    .RESET_B(net155),
    .Q(\line_cache[198][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27955_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01767_),
    .RESET_B(net150),
    .Q(\line_cache[198][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27956_ (.CLK(clknet_leaf_27_clk_i),
    .D(_01768_),
    .RESET_B(net155),
    .Q(\line_cache[198][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27957_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01769_),
    .RESET_B(net149),
    .Q(\line_cache[198][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27958_ (.CLK(clknet_leaf_22_clk_i),
    .D(_01770_),
    .RESET_B(net155),
    .Q(\line_cache[198][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27959_ (.CLK(clknet_leaf_16_clk_i),
    .D(_01771_),
    .RESET_B(net147),
    .Q(\line_cache[199][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27960_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01772_),
    .RESET_B(net147),
    .Q(\line_cache[199][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27961_ (.CLK(clknet_leaf_15_clk_i),
    .D(_01773_),
    .RESET_B(net149),
    .Q(\line_cache[199][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27962_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01774_),
    .RESET_B(net149),
    .Q(\line_cache[199][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27963_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01775_),
    .RESET_B(net149),
    .Q(\line_cache[199][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27964_ (.CLK(clknet_leaf_15_clk_i),
    .D(_01776_),
    .RESET_B(net147),
    .Q(\line_cache[199][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27965_ (.CLK(clknet_leaf_15_clk_i),
    .D(_01777_),
    .RESET_B(net147),
    .Q(\line_cache[199][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27966_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01778_),
    .RESET_B(net149),
    .Q(\line_cache[199][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27967_ (.CLK(clknet_leaf_16_clk_i),
    .D(_01779_),
    .RESET_B(net147),
    .Q(\line_cache[200][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27968_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01780_),
    .RESET_B(net147),
    .Q(\line_cache[200][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27969_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01781_),
    .RESET_B(net147),
    .Q(\line_cache[200][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27970_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01782_),
    .RESET_B(net149),
    .Q(\line_cache[200][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27971_ (.CLK(clknet_leaf_14_clk_i),
    .D(_01783_),
    .RESET_B(net149),
    .Q(\line_cache[200][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27972_ (.CLK(clknet_leaf_16_clk_i),
    .D(_01784_),
    .RESET_B(net147),
    .Q(\line_cache[200][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27973_ (.CLK(clknet_leaf_15_clk_i),
    .D(_01785_),
    .RESET_B(net147),
    .Q(\line_cache[200][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27974_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01786_),
    .RESET_B(net149),
    .Q(\line_cache[200][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27975_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01787_),
    .RESET_B(net148),
    .Q(\line_cache[201][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27976_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01788_),
    .RESET_B(net148),
    .Q(\line_cache[201][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27977_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01789_),
    .RESET_B(net148),
    .Q(\line_cache[201][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27978_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01790_),
    .RESET_B(net149),
    .Q(\line_cache[201][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27979_ (.CLK(clknet_leaf_21_clk_i),
    .D(_01791_),
    .RESET_B(net149),
    .Q(\line_cache[201][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27980_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01792_),
    .RESET_B(net148),
    .Q(\line_cache[201][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27981_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01793_),
    .RESET_B(net148),
    .Q(\line_cache[201][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27982_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01794_),
    .RESET_B(net149),
    .Q(\line_cache[201][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27983_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01795_),
    .RESET_B(net148),
    .Q(\line_cache[202][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27984_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01796_),
    .RESET_B(net148),
    .Q(\line_cache[202][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27985_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01797_),
    .RESET_B(net149),
    .Q(\line_cache[202][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27986_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01798_),
    .RESET_B(net149),
    .Q(\line_cache[202][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27987_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01799_),
    .RESET_B(net149),
    .Q(\line_cache[202][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27988_ (.CLK(clknet_leaf_17_clk_i),
    .D(_01800_),
    .RESET_B(net148),
    .Q(\line_cache[202][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27989_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01801_),
    .RESET_B(net148),
    .Q(\line_cache[202][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27990_ (.CLK(clknet_leaf_20_clk_i),
    .D(_01802_),
    .RESET_B(net150),
    .Q(\line_cache[202][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27991_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01803_),
    .RESET_B(net148),
    .Q(\line_cache[203][0] ));
 sky130_fd_sc_hd__dfrtp_1 _27992_ (.CLK(clknet_leaf_18_clk_i),
    .D(_01804_),
    .RESET_B(net148),
    .Q(\line_cache[203][1] ));
 sky130_fd_sc_hd__dfrtp_1 _27993_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01805_),
    .RESET_B(net156),
    .Q(\line_cache[203][2] ));
 sky130_fd_sc_hd__dfrtp_1 _27994_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01806_),
    .RESET_B(net157),
    .Q(\line_cache[203][3] ));
 sky130_fd_sc_hd__dfrtp_1 _27995_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01807_),
    .RESET_B(net150),
    .Q(\line_cache[203][4] ));
 sky130_fd_sc_hd__dfrtp_1 _27996_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01808_),
    .RESET_B(net148),
    .Q(\line_cache[203][5] ));
 sky130_fd_sc_hd__dfrtp_1 _27997_ (.CLK(clknet_leaf_19_clk_i),
    .D(_01809_),
    .RESET_B(net150),
    .Q(\line_cache[203][6] ));
 sky130_fd_sc_hd__dfrtp_1 _27998_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01810_),
    .RESET_B(net157),
    .Q(\line_cache[203][7] ));
 sky130_fd_sc_hd__dfrtp_1 _27999_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01811_),
    .RESET_B(net188),
    .Q(\line_cache[204][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28000_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01812_),
    .RESET_B(net186),
    .Q(\line_cache[204][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28001_ (.CLK(clknet_leaf_36_clk_i),
    .D(_01813_),
    .RESET_B(net157),
    .Q(\line_cache[204][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28002_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01814_),
    .RESET_B(net188),
    .Q(\line_cache[204][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28003_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01815_),
    .RESET_B(net188),
    .Q(\line_cache[204][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28004_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01816_),
    .RESET_B(net188),
    .Q(\line_cache[204][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28005_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01817_),
    .RESET_B(net157),
    .Q(\line_cache[204][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28006_ (.CLK(clknet_leaf_24_clk_i),
    .D(_01818_),
    .RESET_B(net157),
    .Q(\line_cache[204][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28007_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01819_),
    .RESET_B(net194),
    .Q(\line_cache[205][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28008_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01820_),
    .RESET_B(net194),
    .Q(\line_cache[205][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28009_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01821_),
    .RESET_B(net195),
    .Q(\line_cache[205][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28010_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01822_),
    .RESET_B(net195),
    .Q(\line_cache[205][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28011_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01823_),
    .RESET_B(net194),
    .Q(\line_cache[205][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28012_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01824_),
    .RESET_B(net195),
    .Q(\line_cache[205][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28013_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01825_),
    .RESET_B(net194),
    .Q(\line_cache[205][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28014_ (.CLK(clknet_leaf_25_clk_i),
    .D(_01826_),
    .RESET_B(net157),
    .Q(\line_cache[205][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28015_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01827_),
    .RESET_B(net194),
    .Q(\line_cache[206][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28016_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01828_),
    .RESET_B(net194),
    .Q(\line_cache[206][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28017_ (.CLK(clknet_leaf_59_clk_i),
    .D(_01829_),
    .RESET_B(net195),
    .Q(\line_cache[206][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28018_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01830_),
    .RESET_B(net194),
    .Q(\line_cache[206][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28019_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01831_),
    .RESET_B(net194),
    .Q(\line_cache[206][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28020_ (.CLK(clknet_leaf_60_clk_i),
    .D(_01832_),
    .RESET_B(net195),
    .Q(\line_cache[206][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28021_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01833_),
    .RESET_B(net194),
    .Q(\line_cache[206][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28022_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01834_),
    .RESET_B(net195),
    .Q(\line_cache[206][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28023_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01835_),
    .RESET_B(net188),
    .Q(\line_cache[207][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28024_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01836_),
    .RESET_B(net188),
    .Q(\line_cache[207][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28025_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01837_),
    .RESET_B(net195),
    .Q(\line_cache[207][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28026_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01838_),
    .RESET_B(net195),
    .Q(\line_cache[207][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28027_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01839_),
    .RESET_B(net188),
    .Q(\line_cache[207][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28028_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01840_),
    .RESET_B(net194),
    .Q(\line_cache[207][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28029_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01841_),
    .RESET_B(net188),
    .Q(\line_cache[207][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28030_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01842_),
    .RESET_B(net195),
    .Q(\line_cache[207][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28031_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01843_),
    .RESET_B(net186),
    .Q(\line_cache[208][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28032_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01844_),
    .RESET_B(net186),
    .Q(\line_cache[208][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28033_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01845_),
    .RESET_B(net186),
    .Q(\line_cache[208][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28034_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01846_),
    .RESET_B(net194),
    .Q(\line_cache[208][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28035_ (.CLK(clknet_leaf_65_clk_i),
    .D(_01847_),
    .RESET_B(net188),
    .Q(\line_cache[208][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28036_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01848_),
    .RESET_B(net195),
    .Q(\line_cache[208][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28037_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01849_),
    .RESET_B(net188),
    .Q(\line_cache[208][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28038_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01850_),
    .RESET_B(net194),
    .Q(\line_cache[208][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28039_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01851_),
    .RESET_B(net186),
    .Q(\line_cache[209][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28040_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01852_),
    .RESET_B(net188),
    .Q(\line_cache[209][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28041_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01853_),
    .RESET_B(net188),
    .Q(\line_cache[209][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28042_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01854_),
    .RESET_B(net194),
    .Q(\line_cache[209][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28043_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01855_),
    .RESET_B(net186),
    .Q(\line_cache[209][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28044_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01856_),
    .RESET_B(net194),
    .Q(\line_cache[209][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28045_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01857_),
    .RESET_B(net188),
    .Q(\line_cache[209][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28046_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01858_),
    .RESET_B(net194),
    .Q(\line_cache[209][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28047_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01859_),
    .RESET_B(net186),
    .Q(\line_cache[210][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28048_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01860_),
    .RESET_B(net186),
    .Q(\line_cache[210][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28049_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01861_),
    .RESET_B(net186),
    .Q(\line_cache[210][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28050_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01862_),
    .RESET_B(net197),
    .Q(\line_cache[210][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28051_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01863_),
    .RESET_B(net186),
    .Q(\line_cache[210][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28052_ (.CLK(clknet_leaf_61_clk_i),
    .D(_01864_),
    .RESET_B(net194),
    .Q(\line_cache[210][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28053_ (.CLK(clknet_leaf_66_clk_i),
    .D(_01865_),
    .RESET_B(net188),
    .Q(\line_cache[210][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28054_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01866_),
    .RESET_B(net197),
    .Q(\line_cache[210][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28055_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01867_),
    .RESET_B(net186),
    .Q(\line_cache[211][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28056_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01868_),
    .RESET_B(net186),
    .Q(\line_cache[211][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28057_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01869_),
    .RESET_B(net186),
    .Q(\line_cache[211][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28058_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01870_),
    .RESET_B(net186),
    .Q(\line_cache[211][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28059_ (.CLK(clknet_leaf_67_clk_i),
    .D(_01871_),
    .RESET_B(net186),
    .Q(\line_cache[211][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28060_ (.CLK(clknet_leaf_64_clk_i),
    .D(_01872_),
    .RESET_B(net188),
    .Q(\line_cache[211][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28061_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01873_),
    .RESET_B(net188),
    .Q(\line_cache[211][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28062_ (.CLK(clknet_leaf_63_clk_i),
    .D(_01874_),
    .RESET_B(net189),
    .Q(\line_cache[211][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28063_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01875_),
    .RESET_B(net187),
    .Q(\line_cache[212][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28064_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01876_),
    .RESET_B(net187),
    .Q(\line_cache[212][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28065_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01877_),
    .RESET_B(net187),
    .Q(\line_cache[212][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28066_ (.CLK(clknet_leaf_68_clk_i),
    .D(_01878_),
    .RESET_B(net187),
    .Q(\line_cache[212][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28067_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01879_),
    .RESET_B(net187),
    .Q(\line_cache[212][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28068_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01880_),
    .RESET_B(net189),
    .Q(\line_cache[212][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28069_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01881_),
    .RESET_B(net189),
    .Q(\line_cache[212][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28070_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01882_),
    .RESET_B(net197),
    .Q(\line_cache[212][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28071_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01883_),
    .RESET_B(net187),
    .Q(\line_cache[213][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28072_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01884_),
    .RESET_B(net190),
    .Q(\line_cache[213][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28073_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01885_),
    .RESET_B(net190),
    .Q(\line_cache[213][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28074_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01886_),
    .RESET_B(net187),
    .Q(\line_cache[213][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28075_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01887_),
    .RESET_B(net187),
    .Q(\line_cache[213][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28076_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01888_),
    .RESET_B(net189),
    .Q(\line_cache[213][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28077_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01889_),
    .RESET_B(net189),
    .Q(\line_cache[213][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28078_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01890_),
    .RESET_B(net189),
    .Q(\line_cache[213][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28079_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01891_),
    .RESET_B(net190),
    .Q(\line_cache[214][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28080_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01892_),
    .RESET_B(net190),
    .Q(\line_cache[214][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28081_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01893_),
    .RESET_B(net190),
    .Q(\line_cache[214][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28082_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01894_),
    .RESET_B(net190),
    .Q(\line_cache[214][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28083_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01895_),
    .RESET_B(net187),
    .Q(\line_cache[214][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28084_ (.CLK(clknet_leaf_69_clk_i),
    .D(_01896_),
    .RESET_B(net189),
    .Q(\line_cache[214][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28085_ (.CLK(clknet_leaf_70_clk_i),
    .D(_01897_),
    .RESET_B(net189),
    .Q(\line_cache[214][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28086_ (.CLK(clknet_leaf_63_clk_i),
    .D(_01898_),
    .RESET_B(net189),
    .Q(\line_cache[214][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28087_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01899_),
    .RESET_B(net192),
    .Q(\line_cache[215][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28088_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01900_),
    .RESET_B(net190),
    .Q(\line_cache[215][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28089_ (.CLK(clknet_leaf_72_clk_i),
    .D(_01901_),
    .RESET_B(net190),
    .Q(\line_cache[215][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28090_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01902_),
    .RESET_B(net192),
    .Q(\line_cache[215][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28091_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01903_),
    .RESET_B(net192),
    .Q(\line_cache[215][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28092_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01904_),
    .RESET_B(net192),
    .Q(\line_cache[215][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28093_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01905_),
    .RESET_B(net192),
    .Q(\line_cache[215][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28094_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01906_),
    .RESET_B(net192),
    .Q(\line_cache[215][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28095_ (.CLK(clknet_leaf_71_clk_i),
    .D(_01907_),
    .RESET_B(net192),
    .Q(\line_cache[216][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28096_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01908_),
    .RESET_B(net192),
    .Q(\line_cache[216][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28097_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01909_),
    .RESET_B(net192),
    .Q(\line_cache[216][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28098_ (.CLK(clknet_leaf_78_clk_i),
    .D(_01910_),
    .RESET_B(net197),
    .Q(\line_cache[216][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28099_ (.CLK(clknet_leaf_78_clk_i),
    .D(_01911_),
    .RESET_B(net198),
    .Q(\line_cache[216][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28100_ (.CLK(clknet_leaf_77_clk_i),
    .D(_01912_),
    .RESET_B(net192),
    .Q(\line_cache[216][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28101_ (.CLK(clknet_leaf_78_clk_i),
    .D(_01913_),
    .RESET_B(net198),
    .Q(\line_cache[216][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28102_ (.CLK(clknet_leaf_76_clk_i),
    .D(_01914_),
    .RESET_B(net198),
    .Q(\line_cache[216][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28103_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01915_),
    .RESET_B(net198),
    .Q(\line_cache[217][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28104_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01916_),
    .RESET_B(net198),
    .Q(\line_cache[217][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28105_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01917_),
    .RESET_B(net197),
    .Q(\line_cache[217][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28106_ (.CLK(clknet_leaf_63_clk_i),
    .D(_01918_),
    .RESET_B(net197),
    .Q(\line_cache[217][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28107_ (.CLK(clknet_leaf_56_clk_i),
    .D(_01919_),
    .RESET_B(net198),
    .Q(\line_cache[217][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28108_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01920_),
    .RESET_B(net198),
    .Q(\line_cache[217][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28109_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01921_),
    .RESET_B(net201),
    .Q(\line_cache[217][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28110_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01922_),
    .RESET_B(net201),
    .Q(\line_cache[217][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28111_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01923_),
    .RESET_B(net199),
    .Q(\line_cache[218][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28112_ (.CLK(clknet_leaf_78_clk_i),
    .D(_01924_),
    .RESET_B(net198),
    .Q(\line_cache[218][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28113_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01925_),
    .RESET_B(net195),
    .Q(\line_cache[218][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28114_ (.CLK(clknet_leaf_62_clk_i),
    .D(_01926_),
    .RESET_B(net197),
    .Q(\line_cache[218][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28115_ (.CLK(clknet_leaf_78_clk_i),
    .D(_01927_),
    .RESET_B(net198),
    .Q(\line_cache[218][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28116_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01928_),
    .RESET_B(net201),
    .Q(\line_cache[218][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28117_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01929_),
    .RESET_B(net201),
    .Q(\line_cache[218][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28118_ (.CLK(clknet_leaf_78_clk_i),
    .D(_01930_),
    .RESET_B(net198),
    .Q(\line_cache[218][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28119_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01931_),
    .RESET_B(net195),
    .Q(\line_cache[219][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28120_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01932_),
    .RESET_B(net199),
    .Q(\line_cache[219][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28121_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01933_),
    .RESET_B(net199),
    .Q(\line_cache[219][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28122_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01934_),
    .RESET_B(net199),
    .Q(\line_cache[219][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28123_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01935_),
    .RESET_B(net199),
    .Q(\line_cache[219][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28124_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01936_),
    .RESET_B(net200),
    .Q(\line_cache[219][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28125_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01937_),
    .RESET_B(net200),
    .Q(\line_cache[219][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28126_ (.CLK(clknet_leaf_79_clk_i),
    .D(_01938_),
    .RESET_B(net201),
    .Q(\line_cache[219][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28127_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01939_),
    .RESET_B(net199),
    .Q(\line_cache[220][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28128_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01940_),
    .RESET_B(net199),
    .Q(\line_cache[220][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28129_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01941_),
    .RESET_B(net200),
    .Q(\line_cache[220][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28130_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01942_),
    .RESET_B(net199),
    .Q(\line_cache[220][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28131_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01943_),
    .RESET_B(net199),
    .Q(\line_cache[220][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28132_ (.CLK(clknet_leaf_80_clk_i),
    .D(_01944_),
    .RESET_B(net200),
    .Q(\line_cache[220][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28133_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01945_),
    .RESET_B(net200),
    .Q(\line_cache[220][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28134_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01946_),
    .RESET_B(net200),
    .Q(\line_cache[220][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28135_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01947_),
    .RESET_B(net199),
    .Q(\line_cache[221][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28136_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01948_),
    .RESET_B(net196),
    .Q(\line_cache[221][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28137_ (.CLK(clknet_leaf_55_clk_i),
    .D(_01949_),
    .RESET_B(net199),
    .Q(\line_cache[221][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28138_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01950_),
    .RESET_B(net218),
    .Q(\line_cache[221][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28139_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01951_),
    .RESET_B(net218),
    .Q(\line_cache[221][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28140_ (.CLK(clknet_leaf_54_clk_i),
    .D(_01952_),
    .RESET_B(net199),
    .Q(\line_cache[221][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28141_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01953_),
    .RESET_B(net218),
    .Q(\line_cache[221][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28142_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01954_),
    .RESET_B(net221),
    .Q(\line_cache[221][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28143_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01955_),
    .RESET_B(net199),
    .Q(\line_cache[222][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28144_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01956_),
    .RESET_B(net196),
    .Q(\line_cache[222][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28145_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01957_),
    .RESET_B(net199),
    .Q(\line_cache[222][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28146_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01958_),
    .RESET_B(net218),
    .Q(\line_cache[222][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28147_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01959_),
    .RESET_B(net218),
    .Q(\line_cache[222][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28148_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01960_),
    .RESET_B(net200),
    .Q(\line_cache[222][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28149_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01961_),
    .RESET_B(net221),
    .Q(\line_cache[222][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28150_ (.CLK(clknet_leaf_53_clk_i),
    .D(_01962_),
    .RESET_B(net221),
    .Q(\line_cache[222][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28151_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01963_),
    .RESET_B(net196),
    .Q(\line_cache[223][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28152_ (.CLK(clknet_leaf_52_clk_i),
    .D(_01964_),
    .RESET_B(net218),
    .Q(\line_cache[223][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28153_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01965_),
    .RESET_B(net215),
    .Q(\line_cache[223][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28154_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01966_),
    .RESET_B(net218),
    .Q(\line_cache[223][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28155_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01967_),
    .RESET_B(net218),
    .Q(\line_cache[223][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28156_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01968_),
    .RESET_B(net219),
    .Q(\line_cache[223][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28157_ (.CLK(clknet_leaf_129_clk_i),
    .D(_01969_),
    .RESET_B(net220),
    .Q(\line_cache[223][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28158_ (.CLK(clknet_leaf_131_clk_i),
    .D(_01970_),
    .RESET_B(net220),
    .Q(\line_cache[223][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28159_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01971_),
    .RESET_B(net196),
    .Q(\line_cache[224][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28160_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01972_),
    .RESET_B(net215),
    .Q(\line_cache[224][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28161_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01973_),
    .RESET_B(net196),
    .Q(\line_cache[224][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28162_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01974_),
    .RESET_B(net218),
    .Q(\line_cache[224][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28163_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01975_),
    .RESET_B(net219),
    .Q(\line_cache[224][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28164_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01976_),
    .RESET_B(net219),
    .Q(\line_cache[224][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28165_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01977_),
    .RESET_B(net219),
    .Q(\line_cache[224][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28166_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01978_),
    .RESET_B(net219),
    .Q(\line_cache[224][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28167_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01979_),
    .RESET_B(net196),
    .Q(\line_cache[225][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28168_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01980_),
    .RESET_B(net215),
    .Q(\line_cache[225][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28169_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01981_),
    .RESET_B(net196),
    .Q(\line_cache[225][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28170_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01982_),
    .RESET_B(net217),
    .Q(\line_cache[225][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28171_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01983_),
    .RESET_B(net218),
    .Q(\line_cache[225][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28172_ (.CLK(clknet_leaf_51_clk_i),
    .D(_01984_),
    .RESET_B(net219),
    .Q(\line_cache[225][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28173_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01985_),
    .RESET_B(net216),
    .Q(\line_cache[225][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28174_ (.CLK(clknet_leaf_50_clk_i),
    .D(_01986_),
    .RESET_B(net219),
    .Q(\line_cache[225][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28175_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01987_),
    .RESET_B(net196),
    .Q(\line_cache[226][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28176_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01988_),
    .RESET_B(net217),
    .Q(\line_cache[226][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28177_ (.CLK(clknet_leaf_57_clk_i),
    .D(_01989_),
    .RESET_B(net196),
    .Q(\line_cache[226][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28178_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01990_),
    .RESET_B(net217),
    .Q(\line_cache[226][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28179_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01991_),
    .RESET_B(net217),
    .Q(\line_cache[226][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28180_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01992_),
    .RESET_B(net216),
    .Q(\line_cache[226][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28181_ (.CLK(clknet_leaf_44_clk_i),
    .D(_01993_),
    .RESET_B(net216),
    .Q(\line_cache[226][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28182_ (.CLK(clknet_leaf_49_clk_i),
    .D(_01994_),
    .RESET_B(net216),
    .Q(\line_cache[226][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28183_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01995_),
    .RESET_B(net195),
    .Q(\line_cache[227][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28184_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01996_),
    .RESET_B(net215),
    .Q(\line_cache[227][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28185_ (.CLK(clknet_leaf_58_clk_i),
    .D(_01997_),
    .RESET_B(net196),
    .Q(\line_cache[227][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28186_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01998_),
    .RESET_B(net215),
    .Q(\line_cache[227][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28187_ (.CLK(clknet_leaf_48_clk_i),
    .D(_01999_),
    .RESET_B(net215),
    .Q(\line_cache[227][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28188_ (.CLK(clknet_leaf_48_clk_i),
    .D(_02000_),
    .RESET_B(net215),
    .Q(\line_cache[227][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28189_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02001_),
    .RESET_B(net216),
    .Q(\line_cache[227][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28190_ (.CLK(clknet_leaf_45_clk_i),
    .D(_02002_),
    .RESET_B(net216),
    .Q(\line_cache[227][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28191_ (.CLK(clknet_leaf_58_clk_i),
    .D(_02003_),
    .RESET_B(net195),
    .Q(\line_cache[228][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28192_ (.CLK(clknet_leaf_58_clk_i),
    .D(_02004_),
    .RESET_B(net195),
    .Q(\line_cache[228][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28193_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02005_),
    .RESET_B(net216),
    .Q(\line_cache[228][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28194_ (.CLK(clknet_leaf_48_clk_i),
    .D(_02006_),
    .RESET_B(net215),
    .Q(\line_cache[228][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28195_ (.CLK(clknet_leaf_48_clk_i),
    .D(_02007_),
    .RESET_B(net215),
    .Q(\line_cache[228][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28196_ (.CLK(clknet_leaf_45_clk_i),
    .D(_02008_),
    .RESET_B(net216),
    .Q(\line_cache[228][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28197_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02009_),
    .RESET_B(net216),
    .Q(\line_cache[228][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28198_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02010_),
    .RESET_B(net216),
    .Q(\line_cache[228][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28199_ (.CLK(clknet_leaf_59_clk_i),
    .D(_02011_),
    .RESET_B(net195),
    .Q(\line_cache[229][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28200_ (.CLK(clknet_leaf_48_clk_i),
    .D(_02012_),
    .RESET_B(net215),
    .Q(\line_cache[229][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28201_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02013_),
    .RESET_B(net179),
    .Q(\line_cache[229][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28202_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02014_),
    .RESET_B(net215),
    .Q(\line_cache[229][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28203_ (.CLK(clknet_leaf_36_clk_i),
    .D(_02015_),
    .RESET_B(net178),
    .Q(\line_cache[229][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28204_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02016_),
    .RESET_B(net215),
    .Q(\line_cache[229][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28205_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02017_),
    .RESET_B(net215),
    .Q(\line_cache[229][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28206_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02018_),
    .RESET_B(net179),
    .Q(\line_cache[229][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28207_ (.CLK(clknet_leaf_25_clk_i),
    .D(_02019_),
    .RESET_B(net178),
    .Q(\line_cache[230][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28208_ (.CLK(clknet_leaf_48_clk_i),
    .D(_02020_),
    .RESET_B(net215),
    .Q(\line_cache[230][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28209_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02021_),
    .RESET_B(net179),
    .Q(\line_cache[230][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28210_ (.CLK(clknet_leaf_36_clk_i),
    .D(_02022_),
    .RESET_B(net178),
    .Q(\line_cache[230][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28211_ (.CLK(clknet_leaf_36_clk_i),
    .D(_02023_),
    .RESET_B(net178),
    .Q(\line_cache[230][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28212_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02024_),
    .RESET_B(net215),
    .Q(\line_cache[230][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28213_ (.CLK(clknet_leaf_47_clk_i),
    .D(_02025_),
    .RESET_B(net215),
    .Q(\line_cache[230][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28214_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02026_),
    .RESET_B(net216),
    .Q(\line_cache[230][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28215_ (.CLK(clknet_leaf_36_clk_i),
    .D(_02027_),
    .RESET_B(net180),
    .Q(\line_cache[231][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28216_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02028_),
    .RESET_B(net178),
    .Q(\line_cache[231][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28217_ (.CLK(clknet_leaf_36_clk_i),
    .D(_02029_),
    .RESET_B(net180),
    .Q(\line_cache[231][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28218_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02030_),
    .RESET_B(net178),
    .Q(\line_cache[231][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28219_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02031_),
    .RESET_B(net178),
    .Q(\line_cache[231][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28220_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02032_),
    .RESET_B(net178),
    .Q(\line_cache[231][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28221_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02033_),
    .RESET_B(net180),
    .Q(\line_cache[231][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28222_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02034_),
    .RESET_B(net178),
    .Q(\line_cache[231][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28223_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02035_),
    .RESET_B(net180),
    .Q(\line_cache[232][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28224_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02036_),
    .RESET_B(net178),
    .Q(\line_cache[232][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28225_ (.CLK(clknet_leaf_36_clk_i),
    .D(_02037_),
    .RESET_B(net180),
    .Q(\line_cache[232][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28226_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02038_),
    .RESET_B(net178),
    .Q(\line_cache[232][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28227_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02039_),
    .RESET_B(net175),
    .Q(\line_cache[232][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28228_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02040_),
    .RESET_B(net175),
    .Q(\line_cache[232][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28229_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02041_),
    .RESET_B(net179),
    .Q(\line_cache[232][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28230_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02042_),
    .RESET_B(net178),
    .Q(\line_cache[232][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28231_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02043_),
    .RESET_B(net179),
    .Q(\line_cache[233][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28232_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02044_),
    .RESET_B(net178),
    .Q(\line_cache[233][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28233_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02045_),
    .RESET_B(net179),
    .Q(\line_cache[233][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28234_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02046_),
    .RESET_B(net178),
    .Q(\line_cache[233][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28235_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02047_),
    .RESET_B(net176),
    .Q(\line_cache[233][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28236_ (.CLK(clknet_leaf_33_clk_i),
    .D(_02048_),
    .RESET_B(net176),
    .Q(\line_cache[233][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28237_ (.CLK(clknet_leaf_38_clk_i),
    .D(_02049_),
    .RESET_B(net179),
    .Q(\line_cache[233][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28238_ (.CLK(clknet_leaf_33_clk_i),
    .D(_02050_),
    .RESET_B(net179),
    .Q(\line_cache[233][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28239_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02051_),
    .RESET_B(net179),
    .Q(\line_cache[234][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28240_ (.CLK(clknet_leaf_38_clk_i),
    .D(_02052_),
    .RESET_B(net179),
    .Q(\line_cache[234][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28241_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02053_),
    .RESET_B(net180),
    .Q(\line_cache[234][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28242_ (.CLK(clknet_leaf_33_clk_i),
    .D(_02054_),
    .RESET_B(net179),
    .Q(\line_cache[234][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28243_ (.CLK(clknet_leaf_39_clk_i),
    .D(_02055_),
    .RESET_B(net179),
    .Q(\line_cache[234][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28244_ (.CLK(clknet_leaf_34_clk_i),
    .D(_02056_),
    .RESET_B(net179),
    .Q(\line_cache[234][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28245_ (.CLK(clknet_leaf_38_clk_i),
    .D(_02057_),
    .RESET_B(net179),
    .Q(\line_cache[234][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28246_ (.CLK(clknet_leaf_38_clk_i),
    .D(_02058_),
    .RESET_B(net179),
    .Q(\line_cache[234][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28247_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02059_),
    .RESET_B(net180),
    .Q(\line_cache[235][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28248_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02060_),
    .RESET_B(net180),
    .Q(\line_cache[235][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28249_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02061_),
    .RESET_B(net183),
    .Q(\line_cache[235][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28250_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02062_),
    .RESET_B(net183),
    .Q(\line_cache[235][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28251_ (.CLK(clknet_leaf_39_clk_i),
    .D(_02063_),
    .RESET_B(net183),
    .Q(\line_cache[235][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28252_ (.CLK(clknet_leaf_38_clk_i),
    .D(_02064_),
    .RESET_B(net183),
    .Q(\line_cache[235][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28253_ (.CLK(clknet_leaf_38_clk_i),
    .D(_02065_),
    .RESET_B(net183),
    .Q(\line_cache[235][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28254_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02066_),
    .RESET_B(net183),
    .Q(\line_cache[235][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28255_ (.CLK(clknet_leaf_37_clk_i),
    .D(_02067_),
    .RESET_B(net180),
    .Q(\line_cache[236][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28256_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02068_),
    .RESET_B(net180),
    .Q(\line_cache[236][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28257_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02069_),
    .RESET_B(net222),
    .Q(\line_cache[236][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28258_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02070_),
    .RESET_B(net183),
    .Q(\line_cache[236][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28259_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02071_),
    .RESET_B(net183),
    .Q(\line_cache[236][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28260_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02072_),
    .RESET_B(net183),
    .Q(\line_cache[236][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28261_ (.CLK(clknet_leaf_46_clk_i),
    .D(_02073_),
    .RESET_B(net216),
    .Q(\line_cache[236][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28262_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02074_),
    .RESET_B(net183),
    .Q(\line_cache[236][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28263_ (.CLK(clknet_leaf_45_clk_i),
    .D(_02075_),
    .RESET_B(net216),
    .Q(\line_cache[237][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28264_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02076_),
    .RESET_B(net216),
    .Q(\line_cache[237][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28265_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02077_),
    .RESET_B(net222),
    .Q(\line_cache[237][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28266_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02078_),
    .RESET_B(net222),
    .Q(\line_cache[237][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28267_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02079_),
    .RESET_B(net222),
    .Q(\line_cache[237][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28268_ (.CLK(clknet_leaf_45_clk_i),
    .D(_02080_),
    .RESET_B(net222),
    .Q(\line_cache[237][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28269_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02081_),
    .RESET_B(net222),
    .Q(\line_cache[237][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28270_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02082_),
    .RESET_B(net222),
    .Q(\line_cache[237][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28271_ (.CLK(clknet_leaf_45_clk_i),
    .D(_02083_),
    .RESET_B(net216),
    .Q(\line_cache[238][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28272_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02084_),
    .RESET_B(net217),
    .Q(\line_cache[238][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28273_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02085_),
    .RESET_B(net222),
    .Q(\line_cache[238][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28274_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02086_),
    .RESET_B(net222),
    .Q(\line_cache[238][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28275_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02087_),
    .RESET_B(net222),
    .Q(\line_cache[238][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28276_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02088_),
    .RESET_B(net222),
    .Q(\line_cache[238][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28277_ (.CLK(clknet_leaf_45_clk_i),
    .D(_02089_),
    .RESET_B(net216),
    .Q(\line_cache[238][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28278_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02090_),
    .RESET_B(net222),
    .Q(\line_cache[238][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28279_ (.CLK(clknet_leaf_50_clk_i),
    .D(_02091_),
    .RESET_B(net217),
    .Q(\line_cache[239][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28280_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02092_),
    .RESET_B(net217),
    .Q(\line_cache[239][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28281_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02093_),
    .RESET_B(net222),
    .Q(\line_cache[239][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28282_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02094_),
    .RESET_B(net222),
    .Q(\line_cache[239][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28283_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02095_),
    .RESET_B(net222),
    .Q(\line_cache[239][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28284_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02096_),
    .RESET_B(net222),
    .Q(\line_cache[239][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28285_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02097_),
    .RESET_B(net217),
    .Q(\line_cache[239][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28286_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02098_),
    .RESET_B(net224),
    .Q(\line_cache[239][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28287_ (.CLK(clknet_leaf_50_clk_i),
    .D(_02099_),
    .RESET_B(net219),
    .Q(\line_cache[240][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28288_ (.CLK(clknet_leaf_50_clk_i),
    .D(_02100_),
    .RESET_B(net219),
    .Q(\line_cache[240][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28289_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02101_),
    .RESET_B(net223),
    .Q(\line_cache[240][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28290_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02102_),
    .RESET_B(net223),
    .Q(\line_cache[240][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28291_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02103_),
    .RESET_B(net224),
    .Q(\line_cache[240][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28292_ (.CLK(clknet_leaf_44_clk_i),
    .D(_02104_),
    .RESET_B(net224),
    .Q(\line_cache[240][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28293_ (.CLK(clknet_leaf_50_clk_i),
    .D(_02105_),
    .RESET_B(net217),
    .Q(\line_cache[240][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28294_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02106_),
    .RESET_B(net226),
    .Q(\line_cache[240][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28295_ (.CLK(clknet_leaf_131_clk_i),
    .D(_02107_),
    .RESET_B(net219),
    .Q(\line_cache[241][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28296_ (.CLK(clknet_leaf_131_clk_i),
    .D(_02108_),
    .RESET_B(net219),
    .Q(\line_cache[241][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28297_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02109_),
    .RESET_B(net225),
    .Q(\line_cache[241][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28298_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02110_),
    .RESET_B(net225),
    .Q(\line_cache[241][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28299_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02111_),
    .RESET_B(net225),
    .Q(\line_cache[241][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28300_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02112_),
    .RESET_B(net225),
    .Q(\line_cache[241][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28301_ (.CLK(clknet_leaf_130_clk_i),
    .D(_02113_),
    .RESET_B(net220),
    .Q(\line_cache[241][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28302_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02114_),
    .RESET_B(net225),
    .Q(\line_cache[241][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28303_ (.CLK(clknet_leaf_131_clk_i),
    .D(_02115_),
    .RESET_B(net219),
    .Q(\line_cache[242][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28304_ (.CLK(clknet_leaf_131_clk_i),
    .D(_02116_),
    .RESET_B(net219),
    .Q(\line_cache[242][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28305_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02117_),
    .RESET_B(net225),
    .Q(\line_cache[242][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28306_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02118_),
    .RESET_B(net225),
    .Q(\line_cache[242][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28307_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02119_),
    .RESET_B(net225),
    .Q(\line_cache[242][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28308_ (.CLK(clknet_leaf_131_clk_i),
    .D(_02120_),
    .RESET_B(net219),
    .Q(\line_cache[242][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28309_ (.CLK(clknet_leaf_130_clk_i),
    .D(_02121_),
    .RESET_B(net220),
    .Q(\line_cache[242][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28310_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02122_),
    .RESET_B(net225),
    .Q(\line_cache[242][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28311_ (.CLK(clknet_leaf_133_clk_i),
    .D(_02123_),
    .RESET_B(net227),
    .Q(\line_cache[243][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28312_ (.CLK(clknet_leaf_130_clk_i),
    .D(_02124_),
    .RESET_B(net220),
    .Q(\line_cache[243][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28313_ (.CLK(clknet_leaf_133_clk_i),
    .D(_02125_),
    .RESET_B(net227),
    .Q(\line_cache[243][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28314_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02126_),
    .RESET_B(net225),
    .Q(\line_cache[243][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28315_ (.CLK(clknet_leaf_138_clk_i),
    .D(_02127_),
    .RESET_B(net225),
    .Q(\line_cache[243][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28316_ (.CLK(clknet_leaf_132_clk_i),
    .D(_02128_),
    .RESET_B(net227),
    .Q(\line_cache[243][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28317_ (.CLK(clknet_leaf_133_clk_i),
    .D(_02129_),
    .RESET_B(net227),
    .Q(\line_cache[243][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28318_ (.CLK(clknet_leaf_133_clk_i),
    .D(_02130_),
    .RESET_B(net227),
    .Q(\line_cache[243][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28319_ (.CLK(clknet_leaf_133_clk_i),
    .D(_02131_),
    .RESET_B(net227),
    .Q(\line_cache[244][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28320_ (.CLK(clknet_leaf_134_clk_i),
    .D(_02132_),
    .RESET_B(net226),
    .Q(\line_cache[244][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28321_ (.CLK(clknet_leaf_133_clk_i),
    .D(_02133_),
    .RESET_B(net227),
    .Q(\line_cache[244][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28322_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02134_),
    .RESET_B(net226),
    .Q(\line_cache[244][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28323_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02135_),
    .RESET_B(net226),
    .Q(\line_cache[244][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28324_ (.CLK(clknet_leaf_136_clk_i),
    .D(_02136_),
    .RESET_B(net226),
    .Q(\line_cache[244][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28325_ (.CLK(clknet_leaf_135_clk_i),
    .D(_02137_),
    .RESET_B(net226),
    .Q(\line_cache[244][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28326_ (.CLK(clknet_leaf_135_clk_i),
    .D(_02138_),
    .RESET_B(net226),
    .Q(\line_cache[244][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28327_ (.CLK(clknet_leaf_134_clk_i),
    .D(_02139_),
    .RESET_B(net226),
    .Q(\line_cache[245][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28328_ (.CLK(clknet_leaf_135_clk_i),
    .D(_02140_),
    .RESET_B(net226),
    .Q(\line_cache[245][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28329_ (.CLK(clknet_leaf_121_clk_i),
    .D(_02141_),
    .RESET_B(net236),
    .Q(\line_cache[245][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28330_ (.CLK(clknet_leaf_136_clk_i),
    .D(_02142_),
    .RESET_B(net226),
    .Q(\line_cache[245][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28331_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02143_),
    .RESET_B(net226),
    .Q(\line_cache[245][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28332_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02144_),
    .RESET_B(net305),
    .Q(\line_cache[245][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28333_ (.CLK(clknet_leaf_134_clk_i),
    .D(_02145_),
    .RESET_B(net226),
    .Q(\line_cache[245][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28334_ (.CLK(clknet_leaf_135_clk_i),
    .D(_02146_),
    .RESET_B(net305),
    .Q(\line_cache[245][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28335_ (.CLK(clknet_leaf_134_clk_i),
    .D(_02147_),
    .RESET_B(net226),
    .Q(\line_cache[246][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28336_ (.CLK(clknet_leaf_134_clk_i),
    .D(_02148_),
    .RESET_B(net227),
    .Q(\line_cache[246][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28337_ (.CLK(clknet_leaf_122_clk_i),
    .D(_02149_),
    .RESET_B(net236),
    .Q(\line_cache[246][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28338_ (.CLK(clknet_leaf_136_clk_i),
    .D(_02150_),
    .RESET_B(net304),
    .Q(\line_cache[246][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28339_ (.CLK(clknet_leaf_136_clk_i),
    .D(_02151_),
    .RESET_B(net226),
    .Q(\line_cache[246][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28340_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02152_),
    .RESET_B(net304),
    .Q(\line_cache[246][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28341_ (.CLK(clknet_leaf_121_clk_i),
    .D(_02153_),
    .RESET_B(net237),
    .Q(\line_cache[246][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28342_ (.CLK(clknet_leaf_157_clk_i),
    .D(_02154_),
    .RESET_B(net316),
    .Q(\line_cache[246][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28343_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02155_),
    .RESET_B(net305),
    .Q(\line_cache[247][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28344_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02156_),
    .RESET_B(net305),
    .Q(\line_cache[247][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28345_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02157_),
    .RESET_B(net305),
    .Q(\line_cache[247][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28346_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02158_),
    .RESET_B(net304),
    .Q(\line_cache[247][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28347_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02159_),
    .RESET_B(net304),
    .Q(\line_cache[247][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28348_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02160_),
    .RESET_B(net304),
    .Q(\line_cache[247][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28349_ (.CLK(clknet_leaf_146_clk_i),
    .D(_02161_),
    .RESET_B(net305),
    .Q(\line_cache[247][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28350_ (.CLK(clknet_leaf_146_clk_i),
    .D(_02162_),
    .RESET_B(net305),
    .Q(\line_cache[247][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28351_ (.CLK(clknet_leaf_146_clk_i),
    .D(_02163_),
    .RESET_B(net305),
    .Q(\line_cache[248][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28352_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02164_),
    .RESET_B(net305),
    .Q(\line_cache[248][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28353_ (.CLK(clknet_leaf_146_clk_i),
    .D(_02165_),
    .RESET_B(net305),
    .Q(\line_cache[248][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28354_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02166_),
    .RESET_B(net304),
    .Q(\line_cache[248][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28355_ (.CLK(clknet_leaf_144_clk_i),
    .D(_02167_),
    .RESET_B(net304),
    .Q(\line_cache[248][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28356_ (.CLK(clknet_leaf_145_clk_i),
    .D(_02168_),
    .RESET_B(net304),
    .Q(\line_cache[248][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28357_ (.CLK(clknet_leaf_146_clk_i),
    .D(_02169_),
    .RESET_B(net305),
    .Q(\line_cache[248][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28358_ (.CLK(clknet_leaf_144_clk_i),
    .D(_02170_),
    .RESET_B(net304),
    .Q(\line_cache[248][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28359_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02171_),
    .RESET_B(net304),
    .Q(\line_cache[249][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28360_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02172_),
    .RESET_B(net226),
    .Q(\line_cache[249][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28361_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02173_),
    .RESET_B(net223),
    .Q(\line_cache[249][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28362_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02174_),
    .RESET_B(net223),
    .Q(\line_cache[249][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28363_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02175_),
    .RESET_B(net223),
    .Q(\line_cache[249][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28364_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02176_),
    .RESET_B(net301),
    .Q(\line_cache[249][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28365_ (.CLK(clknet_leaf_144_clk_i),
    .D(_02177_),
    .RESET_B(net304),
    .Q(\line_cache[249][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28366_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02178_),
    .RESET_B(net301),
    .Q(\line_cache[249][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28367_ (.CLK(clknet_leaf_144_clk_i),
    .D(_02179_),
    .RESET_B(net304),
    .Q(\line_cache[250][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28368_ (.CLK(clknet_leaf_137_clk_i),
    .D(_02180_),
    .RESET_B(net226),
    .Q(\line_cache[250][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28369_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02181_),
    .RESET_B(net301),
    .Q(\line_cache[250][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28370_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02182_),
    .RESET_B(net224),
    .Q(\line_cache[250][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28371_ (.CLK(clknet_leaf_139_clk_i),
    .D(_02183_),
    .RESET_B(net224),
    .Q(\line_cache[250][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28372_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02184_),
    .RESET_B(net301),
    .Q(\line_cache[250][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28373_ (.CLK(clknet_leaf_144_clk_i),
    .D(_02185_),
    .RESET_B(net304),
    .Q(\line_cache[250][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28374_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02186_),
    .RESET_B(net301),
    .Q(\line_cache[250][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28375_ (.CLK(clknet_leaf_143_clk_i),
    .D(_02187_),
    .RESET_B(net303),
    .Q(\line_cache[251][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28376_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02188_),
    .RESET_B(net303),
    .Q(\line_cache[251][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28377_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02189_),
    .RESET_B(net303),
    .Q(\line_cache[251][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28378_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02190_),
    .RESET_B(net224),
    .Q(\line_cache[251][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28379_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02191_),
    .RESET_B(net224),
    .Q(\line_cache[251][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28380_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02192_),
    .RESET_B(net303),
    .Q(\line_cache[251][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28381_ (.CLK(clknet_leaf_143_clk_i),
    .D(_02193_),
    .RESET_B(net303),
    .Q(\line_cache[251][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28382_ (.CLK(clknet_leaf_143_clk_i),
    .D(_02194_),
    .RESET_B(net303),
    .Q(\line_cache[251][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28383_ (.CLK(clknet_leaf_143_clk_i),
    .D(_02195_),
    .RESET_B(net303),
    .Q(\line_cache[252][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28384_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02196_),
    .RESET_B(net303),
    .Q(\line_cache[252][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28385_ (.CLK(clknet_leaf_141_clk_i),
    .D(_02197_),
    .RESET_B(net301),
    .Q(\line_cache[252][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28386_ (.CLK(clknet_leaf_142_clk_i),
    .D(_02198_),
    .RESET_B(net303),
    .Q(\line_cache[252][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28387_ (.CLK(clknet_leaf_226_clk_i),
    .D(_02199_),
    .RESET_B(net302),
    .Q(\line_cache[252][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28388_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02200_),
    .RESET_B(net301),
    .Q(\line_cache[252][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28389_ (.CLK(clknet_leaf_143_clk_i),
    .D(_02201_),
    .RESET_B(net303),
    .Q(\line_cache[252][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28390_ (.CLK(clknet_leaf_143_clk_i),
    .D(_02202_),
    .RESET_B(net303),
    .Q(\line_cache[252][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28391_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02203_),
    .RESET_B(net302),
    .Q(\line_cache[253][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28392_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02204_),
    .RESET_B(net301),
    .Q(\line_cache[253][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28393_ (.CLK(clknet_leaf_226_clk_i),
    .D(_02205_),
    .RESET_B(net302),
    .Q(\line_cache[253][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28394_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02206_),
    .RESET_B(net302),
    .Q(\line_cache[253][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28395_ (.CLK(clknet_leaf_227_clk_i),
    .D(_02207_),
    .RESET_B(net302),
    .Q(\line_cache[253][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28396_ (.CLK(clknet_leaf_223_clk_i),
    .D(_02208_),
    .RESET_B(net307),
    .Q(\line_cache[253][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28397_ (.CLK(clknet_leaf_226_clk_i),
    .D(_02209_),
    .RESET_B(net307),
    .Q(\line_cache[253][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28398_ (.CLK(clknet_leaf_226_clk_i),
    .D(_02210_),
    .RESET_B(net302),
    .Q(\line_cache[253][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28399_ (.CLK(clknet_leaf_226_clk_i),
    .D(_02211_),
    .RESET_B(net302),
    .Q(\line_cache[254][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28400_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02212_),
    .RESET_B(net302),
    .Q(\line_cache[254][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28401_ (.CLK(clknet_leaf_227_clk_i),
    .D(_02213_),
    .RESET_B(net302),
    .Q(\line_cache[254][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28402_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02214_),
    .RESET_B(net261),
    .Q(\line_cache[254][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28403_ (.CLK(clknet_leaf_227_clk_i),
    .D(_02215_),
    .RESET_B(net302),
    .Q(\line_cache[254][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28404_ (.CLK(clknet_leaf_223_clk_i),
    .D(_02216_),
    .RESET_B(net307),
    .Q(\line_cache[254][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28405_ (.CLK(clknet_leaf_223_clk_i),
    .D(_02217_),
    .RESET_B(net307),
    .Q(\line_cache[254][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28406_ (.CLK(clknet_leaf_226_clk_i),
    .D(_02218_),
    .RESET_B(net302),
    .Q(\line_cache[254][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28407_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02219_),
    .RESET_B(net261),
    .Q(\line_cache[255][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28408_ (.CLK(clknet_leaf_318_clk_i),
    .D(_02220_),
    .RESET_B(net259),
    .Q(\line_cache[255][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28409_ (.CLK(clknet_leaf_317_clk_i),
    .D(_02221_),
    .RESET_B(net259),
    .Q(\line_cache[255][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28410_ (.CLK(clknet_leaf_318_clk_i),
    .D(_02222_),
    .RESET_B(net259),
    .Q(\line_cache[255][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28411_ (.CLK(clknet_leaf_317_clk_i),
    .D(_02223_),
    .RESET_B(net259),
    .Q(\line_cache[255][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28412_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02224_),
    .RESET_B(net261),
    .Q(\line_cache[255][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28413_ (.CLK(clknet_leaf_231_clk_i),
    .D(_02225_),
    .RESET_B(net267),
    .Q(\line_cache[255][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28414_ (.CLK(clknet_leaf_231_clk_i),
    .D(_02226_),
    .RESET_B(net267),
    .Q(\line_cache[255][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28415_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02227_),
    .RESET_B(net181),
    .Q(\line_cache[256][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28416_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02228_),
    .RESET_B(net181),
    .Q(\line_cache[256][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28417_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02229_),
    .RESET_B(net172),
    .Q(\line_cache[256][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28418_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02230_),
    .RESET_B(net181),
    .Q(\line_cache[256][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28419_ (.CLK(clknet_leaf_339_clk_i),
    .D(_02231_),
    .RESET_B(net171),
    .Q(\line_cache[256][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28420_ (.CLK(clknet_leaf_339_clk_i),
    .D(_02232_),
    .RESET_B(net172),
    .Q(\line_cache[256][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28421_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02233_),
    .RESET_B(net248),
    .Q(\line_cache[256][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28422_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02234_),
    .RESET_B(net248),
    .Q(\line_cache[256][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28423_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02235_),
    .RESET_B(net223),
    .Q(\line_cache[257][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28424_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02236_),
    .RESET_B(net223),
    .Q(\line_cache[257][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28425_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02237_),
    .RESET_B(net184),
    .Q(\line_cache[257][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28426_ (.CLK(clknet_leaf_41_clk_i),
    .D(_02238_),
    .RESET_B(net184),
    .Q(\line_cache[257][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28427_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02239_),
    .RESET_B(net223),
    .Q(\line_cache[257][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28428_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02240_),
    .RESET_B(net260),
    .Q(\line_cache[257][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28429_ (.CLK(clknet_leaf_141_clk_i),
    .D(_02241_),
    .RESET_B(net301),
    .Q(\line_cache[257][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28430_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02242_),
    .RESET_B(net301),
    .Q(\line_cache[257][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28431_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02243_),
    .RESET_B(net301),
    .Q(\line_cache[258][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28432_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02244_),
    .RESET_B(net223),
    .Q(\line_cache[258][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28433_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02245_),
    .RESET_B(net184),
    .Q(\line_cache[258][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28434_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02246_),
    .RESET_B(net223),
    .Q(\line_cache[258][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28435_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02247_),
    .RESET_B(net223),
    .Q(\line_cache[258][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28436_ (.CLK(clknet_leaf_41_clk_i),
    .D(_02248_),
    .RESET_B(net184),
    .Q(\line_cache[258][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28437_ (.CLK(clknet_leaf_141_clk_i),
    .D(_02249_),
    .RESET_B(net301),
    .Q(\line_cache[258][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28438_ (.CLK(clknet_leaf_141_clk_i),
    .D(_02250_),
    .RESET_B(net301),
    .Q(\line_cache[258][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28439_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02251_),
    .RESET_B(net223),
    .Q(\line_cache[259][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28440_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02252_),
    .RESET_B(net223),
    .Q(\line_cache[259][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28441_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02253_),
    .RESET_B(net184),
    .Q(\line_cache[259][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28442_ (.CLK(clknet_leaf_43_clk_i),
    .D(_02254_),
    .RESET_B(net184),
    .Q(\line_cache[259][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28443_ (.CLK(clknet_leaf_140_clk_i),
    .D(_02255_),
    .RESET_B(net223),
    .Q(\line_cache[259][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28444_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02256_),
    .RESET_B(net260),
    .Q(\line_cache[259][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28445_ (.CLK(clknet_leaf_141_clk_i),
    .D(_02257_),
    .RESET_B(net301),
    .Q(\line_cache[259][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28446_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02258_),
    .RESET_B(net301),
    .Q(\line_cache[259][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28447_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02259_),
    .RESET_B(net223),
    .Q(\line_cache[260][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28448_ (.CLK(clknet_leaf_42_clk_i),
    .D(_02260_),
    .RESET_B(net223),
    .Q(\line_cache[260][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28449_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02261_),
    .RESET_B(net260),
    .Q(\line_cache[260][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28450_ (.CLK(clknet_leaf_41_clk_i),
    .D(_02262_),
    .RESET_B(net184),
    .Q(\line_cache[260][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28451_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02263_),
    .RESET_B(net301),
    .Q(\line_cache[260][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28452_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02264_),
    .RESET_B(net261),
    .Q(\line_cache[260][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28453_ (.CLK(clknet_leaf_228_clk_i),
    .D(_02265_),
    .RESET_B(net260),
    .Q(\line_cache[260][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28454_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02266_),
    .RESET_B(net260),
    .Q(\line_cache[260][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28455_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02267_),
    .RESET_B(net184),
    .Q(\line_cache[261][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28456_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02268_),
    .RESET_B(net184),
    .Q(\line_cache[261][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28457_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02269_),
    .RESET_B(net184),
    .Q(\line_cache[261][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28458_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02270_),
    .RESET_B(net184),
    .Q(\line_cache[261][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28459_ (.CLK(clknet_leaf_328_clk_i),
    .D(_02271_),
    .RESET_B(net183),
    .Q(\line_cache[261][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28460_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02272_),
    .RESET_B(net260),
    .Q(\line_cache[261][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28461_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02273_),
    .RESET_B(net260),
    .Q(\line_cache[261][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28462_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02274_),
    .RESET_B(net261),
    .Q(\line_cache[261][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28463_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02275_),
    .RESET_B(net184),
    .Q(\line_cache[262][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28464_ (.CLK(clknet_leaf_41_clk_i),
    .D(_02276_),
    .RESET_B(net184),
    .Q(\line_cache[262][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28465_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02277_),
    .RESET_B(net184),
    .Q(\line_cache[262][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28466_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02278_),
    .RESET_B(net185),
    .Q(\line_cache[262][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28467_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02279_),
    .RESET_B(net183),
    .Q(\line_cache[262][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28468_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02280_),
    .RESET_B(net260),
    .Q(\line_cache[262][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28469_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02281_),
    .RESET_B(net261),
    .Q(\line_cache[262][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28470_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02282_),
    .RESET_B(net261),
    .Q(\line_cache[262][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28471_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02283_),
    .RESET_B(net185),
    .Q(\line_cache[263][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28472_ (.CLK(clknet_leaf_41_clk_i),
    .D(_02284_),
    .RESET_B(net185),
    .Q(\line_cache[263][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28473_ (.CLK(clknet_leaf_328_clk_i),
    .D(_02285_),
    .RESET_B(net185),
    .Q(\line_cache[263][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28474_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02286_),
    .RESET_B(net185),
    .Q(\line_cache[263][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28475_ (.CLK(clknet_leaf_328_clk_i),
    .D(_02287_),
    .RESET_B(net185),
    .Q(\line_cache[263][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28476_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02288_),
    .RESET_B(net260),
    .Q(\line_cache[263][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28477_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02289_),
    .RESET_B(net260),
    .Q(\line_cache[263][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28478_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02290_),
    .RESET_B(net261),
    .Q(\line_cache[263][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28479_ (.CLK(clknet_leaf_326_clk_i),
    .D(_02291_),
    .RESET_B(net260),
    .Q(\line_cache[264][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28480_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02292_),
    .RESET_B(net184),
    .Q(\line_cache[264][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28481_ (.CLK(clknet_leaf_40_clk_i),
    .D(_02293_),
    .RESET_B(net183),
    .Q(\line_cache[264][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28482_ (.CLK(clknet_leaf_327_clk_i),
    .D(_02294_),
    .RESET_B(net185),
    .Q(\line_cache[264][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28483_ (.CLK(clknet_leaf_328_clk_i),
    .D(_02295_),
    .RESET_B(net183),
    .Q(\line_cache[264][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28484_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02296_),
    .RESET_B(net260),
    .Q(\line_cache[264][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28485_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02297_),
    .RESET_B(net260),
    .Q(\line_cache[264][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28486_ (.CLK(clknet_leaf_325_clk_i),
    .D(_02298_),
    .RESET_B(net261),
    .Q(\line_cache[264][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28487_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02299_),
    .RESET_B(net261),
    .Q(\line_cache[265][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28488_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02300_),
    .RESET_B(net261),
    .Q(\line_cache[265][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28489_ (.CLK(clknet_leaf_231_clk_i),
    .D(_02301_),
    .RESET_B(net261),
    .Q(\line_cache[265][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28490_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02302_),
    .RESET_B(net259),
    .Q(\line_cache[265][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28491_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02303_),
    .RESET_B(net261),
    .Q(\line_cache[265][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28492_ (.CLK(clknet_leaf_236_clk_i),
    .D(_02304_),
    .RESET_B(net264),
    .Q(\line_cache[265][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28493_ (.CLK(clknet_leaf_235_clk_i),
    .D(_02305_),
    .RESET_B(net265),
    .Q(\line_cache[265][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28494_ (.CLK(clknet_leaf_231_clk_i),
    .D(_02306_),
    .RESET_B(net267),
    .Q(\line_cache[265][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28495_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02307_),
    .RESET_B(net261),
    .Q(\line_cache[266][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28496_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02308_),
    .RESET_B(net261),
    .Q(\line_cache[266][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28497_ (.CLK(clknet_leaf_229_clk_i),
    .D(_02309_),
    .RESET_B(net262),
    .Q(\line_cache[266][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28498_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02310_),
    .RESET_B(net262),
    .Q(\line_cache[266][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28499_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02311_),
    .RESET_B(net262),
    .Q(\line_cache[266][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28500_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02312_),
    .RESET_B(net265),
    .Q(\line_cache[266][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28501_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02313_),
    .RESET_B(net265),
    .Q(\line_cache[266][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28502_ (.CLK(clknet_leaf_231_clk_i),
    .D(_02314_),
    .RESET_B(net267),
    .Q(\line_cache[266][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28503_ (.CLK(clknet_leaf_324_clk_i),
    .D(_02315_),
    .RESET_B(net260),
    .Q(\line_cache[267][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28504_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02316_),
    .RESET_B(net262),
    .Q(\line_cache[267][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28505_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02317_),
    .RESET_B(net262),
    .Q(\line_cache[267][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28506_ (.CLK(clknet_leaf_322_clk_i),
    .D(_02318_),
    .RESET_B(net262),
    .Q(\line_cache[267][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28507_ (.CLK(clknet_leaf_322_clk_i),
    .D(_02319_),
    .RESET_B(net262),
    .Q(\line_cache[267][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28508_ (.CLK(clknet_leaf_318_clk_i),
    .D(_02320_),
    .RESET_B(net264),
    .Q(\line_cache[267][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28509_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02321_),
    .RESET_B(net265),
    .Q(\line_cache[267][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28510_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02322_),
    .RESET_B(net265),
    .Q(\line_cache[267][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28511_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02323_),
    .RESET_B(net260),
    .Q(\line_cache[268][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28512_ (.CLK(clknet_leaf_323_clk_i),
    .D(_02324_),
    .RESET_B(net260),
    .Q(\line_cache[268][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28513_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02325_),
    .RESET_B(net262),
    .Q(\line_cache[268][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28514_ (.CLK(clknet_leaf_322_clk_i),
    .D(_02326_),
    .RESET_B(net258),
    .Q(\line_cache[268][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28515_ (.CLK(clknet_leaf_322_clk_i),
    .D(_02327_),
    .RESET_B(net262),
    .Q(\line_cache[268][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28516_ (.CLK(clknet_leaf_318_clk_i),
    .D(_02328_),
    .RESET_B(net264),
    .Q(\line_cache[268][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28517_ (.CLK(clknet_leaf_318_clk_i),
    .D(_02329_),
    .RESET_B(net264),
    .Q(\line_cache[268][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28518_ (.CLK(clknet_leaf_230_clk_i),
    .D(_02330_),
    .RESET_B(net265),
    .Q(\line_cache[268][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28519_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02331_),
    .RESET_B(net181),
    .Q(\line_cache[269][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28520_ (.CLK(clknet_leaf_329_clk_i),
    .D(_02332_),
    .RESET_B(net181),
    .Q(\line_cache[269][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28521_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02333_),
    .RESET_B(net181),
    .Q(\line_cache[269][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28522_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02334_),
    .RESET_B(net182),
    .Q(\line_cache[269][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28523_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02335_),
    .RESET_B(net182),
    .Q(\line_cache[269][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28524_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02336_),
    .RESET_B(net182),
    .Q(\line_cache[269][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28525_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02337_),
    .RESET_B(net258),
    .Q(\line_cache[269][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28526_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02338_),
    .RESET_B(net258),
    .Q(\line_cache[269][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28527_ (.CLK(clknet_leaf_329_clk_i),
    .D(_02339_),
    .RESET_B(net182),
    .Q(\line_cache[270][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28528_ (.CLK(clknet_leaf_329_clk_i),
    .D(_02340_),
    .RESET_B(net182),
    .Q(\line_cache[270][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28529_ (.CLK(clknet_leaf_329_clk_i),
    .D(_02341_),
    .RESET_B(net258),
    .Q(\line_cache[270][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28530_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02342_),
    .RESET_B(net182),
    .Q(\line_cache[270][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28531_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02343_),
    .RESET_B(net258),
    .Q(\line_cache[270][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28532_ (.CLK(clknet_leaf_330_clk_i),
    .D(_02344_),
    .RESET_B(net182),
    .Q(\line_cache[270][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28533_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02345_),
    .RESET_B(net258),
    .Q(\line_cache[270][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28534_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02346_),
    .RESET_B(net259),
    .Q(\line_cache[270][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28535_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02347_),
    .RESET_B(net259),
    .Q(\line_cache[271][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28536_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02348_),
    .RESET_B(net258),
    .Q(\line_cache[271][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28537_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02349_),
    .RESET_B(net259),
    .Q(\line_cache[271][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28538_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02350_),
    .RESET_B(net258),
    .Q(\line_cache[271][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28539_ (.CLK(clknet_leaf_322_clk_i),
    .D(_02351_),
    .RESET_B(net259),
    .Q(\line_cache[271][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28540_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02352_),
    .RESET_B(net258),
    .Q(\line_cache[271][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28541_ (.CLK(clknet_leaf_322_clk_i),
    .D(_02353_),
    .RESET_B(net259),
    .Q(\line_cache[271][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28542_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02354_),
    .RESET_B(net258),
    .Q(\line_cache[271][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28543_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02355_),
    .RESET_B(net175),
    .Q(\line_cache[272][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28544_ (.CLK(clknet_leaf_28_clk_i),
    .D(_02356_),
    .RESET_B(net154),
    .Q(\line_cache[272][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28545_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02357_),
    .RESET_B(net154),
    .Q(\line_cache[272][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28546_ (.CLK(clknet_leaf_28_clk_i),
    .D(_02358_),
    .RESET_B(net152),
    .Q(\line_cache[272][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28547_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02359_),
    .RESET_B(net175),
    .Q(\line_cache[272][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28548_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02360_),
    .RESET_B(net175),
    .Q(\line_cache[272][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28549_ (.CLK(clknet_leaf_333_clk_i),
    .D(_02361_),
    .RESET_B(net176),
    .Q(\line_cache[272][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28550_ (.CLK(clknet_leaf_333_clk_i),
    .D(_02362_),
    .RESET_B(net176),
    .Q(\line_cache[272][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28551_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02363_),
    .RESET_B(net154),
    .Q(\line_cache[273][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28552_ (.CLK(clknet_leaf_28_clk_i),
    .D(_02364_),
    .RESET_B(net154),
    .Q(\line_cache[273][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28553_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02365_),
    .RESET_B(net154),
    .Q(\line_cache[273][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28554_ (.CLK(clknet_leaf_10_clk_i),
    .D(_02366_),
    .RESET_B(net154),
    .Q(\line_cache[273][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28555_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02367_),
    .RESET_B(net175),
    .Q(\line_cache[273][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28556_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02368_),
    .RESET_B(net175),
    .Q(\line_cache[273][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28557_ (.CLK(clknet_leaf_333_clk_i),
    .D(_02369_),
    .RESET_B(net176),
    .Q(\line_cache[273][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28558_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02370_),
    .RESET_B(net176),
    .Q(\line_cache[273][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28559_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02371_),
    .RESET_B(net153),
    .Q(\line_cache[274][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28560_ (.CLK(clknet_leaf_10_clk_i),
    .D(_02372_),
    .RESET_B(net151),
    .Q(\line_cache[274][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28561_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02373_),
    .RESET_B(net153),
    .Q(\line_cache[274][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28562_ (.CLK(clknet_leaf_10_clk_i),
    .D(_02374_),
    .RESET_B(net151),
    .Q(\line_cache[274][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28563_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02375_),
    .RESET_B(net175),
    .Q(\line_cache[274][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28564_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02376_),
    .RESET_B(net175),
    .Q(\line_cache[274][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28565_ (.CLK(clknet_leaf_333_clk_i),
    .D(_02377_),
    .RESET_B(net176),
    .Q(\line_cache[274][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28566_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02378_),
    .RESET_B(net176),
    .Q(\line_cache[274][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28567_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02379_),
    .RESET_B(net153),
    .Q(\line_cache[275][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28568_ (.CLK(clknet_leaf_10_clk_i),
    .D(_02380_),
    .RESET_B(net151),
    .Q(\line_cache[275][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28569_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02381_),
    .RESET_B(net153),
    .Q(\line_cache[275][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28570_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02382_),
    .RESET_B(net153),
    .Q(\line_cache[275][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28571_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02383_),
    .RESET_B(net175),
    .Q(\line_cache[275][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28572_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02384_),
    .RESET_B(net175),
    .Q(\line_cache[275][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28573_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02385_),
    .RESET_B(net176),
    .Q(\line_cache[275][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28574_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02386_),
    .RESET_B(net176),
    .Q(\line_cache[275][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28575_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02387_),
    .RESET_B(net153),
    .Q(\line_cache[276][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28576_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02388_),
    .RESET_B(net153),
    .Q(\line_cache[276][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28577_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02389_),
    .RESET_B(net153),
    .Q(\line_cache[276][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28578_ (.CLK(clknet_leaf_10_clk_i),
    .D(_02390_),
    .RESET_B(net153),
    .Q(\line_cache[276][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28579_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02391_),
    .RESET_B(net175),
    .Q(\line_cache[276][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28580_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02392_),
    .RESET_B(net175),
    .Q(\line_cache[276][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28581_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02393_),
    .RESET_B(net176),
    .Q(\line_cache[276][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28582_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02394_),
    .RESET_B(net176),
    .Q(\line_cache[276][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28583_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02395_),
    .RESET_B(net143),
    .Q(\line_cache[277][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28584_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02396_),
    .RESET_B(net143),
    .Q(\line_cache[277][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28585_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02397_),
    .RESET_B(net153),
    .Q(\line_cache[277][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28586_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02398_),
    .RESET_B(net143),
    .Q(\line_cache[277][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28587_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02399_),
    .RESET_B(net163),
    .Q(\line_cache[277][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28588_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02400_),
    .RESET_B(net163),
    .Q(\line_cache[277][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28589_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02401_),
    .RESET_B(net164),
    .Q(\line_cache[277][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28590_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02402_),
    .RESET_B(net164),
    .Q(\line_cache[277][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28591_ (.CLK(clknet_leaf_362_clk_i),
    .D(_02403_),
    .RESET_B(net143),
    .Q(\line_cache[278][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28592_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02404_),
    .RESET_B(net143),
    .Q(\line_cache[278][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28593_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02405_),
    .RESET_B(net144),
    .Q(\line_cache[278][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28594_ (.CLK(clknet_leaf_7_clk_i),
    .D(_02406_),
    .RESET_B(net144),
    .Q(\line_cache[278][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28595_ (.CLK(clknet_leaf_361_clk_i),
    .D(_02407_),
    .RESET_B(net163),
    .Q(\line_cache[278][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28596_ (.CLK(clknet_leaf_361_clk_i),
    .D(_02408_),
    .RESET_B(net163),
    .Q(\line_cache[278][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28597_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02409_),
    .RESET_B(net164),
    .Q(\line_cache[278][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28598_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02410_),
    .RESET_B(net165),
    .Q(\line_cache[278][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28599_ (.CLK(clknet_leaf_362_clk_i),
    .D(_02411_),
    .RESET_B(net144),
    .Q(\line_cache[279][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28600_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02412_),
    .RESET_B(net144),
    .Q(\line_cache[279][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28601_ (.CLK(clknet_leaf_8_clk_i),
    .D(_02413_),
    .RESET_B(net144),
    .Q(\line_cache[279][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28602_ (.CLK(clknet_leaf_7_clk_i),
    .D(_02414_),
    .RESET_B(net145),
    .Q(\line_cache[279][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28603_ (.CLK(clknet_leaf_360_clk_i),
    .D(_02415_),
    .RESET_B(net163),
    .Q(\line_cache[279][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28604_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02416_),
    .RESET_B(net163),
    .Q(\line_cache[279][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28605_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02417_),
    .RESET_B(net165),
    .Q(\line_cache[279][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28606_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02418_),
    .RESET_B(net165),
    .Q(\line_cache[279][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28607_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02419_),
    .RESET_B(net143),
    .Q(\line_cache[280][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28608_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02420_),
    .RESET_B(net143),
    .Q(\line_cache[280][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28609_ (.CLK(clknet_leaf_362_clk_i),
    .D(_02421_),
    .RESET_B(net144),
    .Q(\line_cache[280][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28610_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02422_),
    .RESET_B(net143),
    .Q(\line_cache[280][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28611_ (.CLK(clknet_leaf_361_clk_i),
    .D(_02423_),
    .RESET_B(net163),
    .Q(\line_cache[280][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28612_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02424_),
    .RESET_B(net164),
    .Q(\line_cache[280][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28613_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02425_),
    .RESET_B(net164),
    .Q(\line_cache[280][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28614_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02426_),
    .RESET_B(net164),
    .Q(\line_cache[280][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28615_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02427_),
    .RESET_B(net143),
    .Q(\line_cache[281][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28616_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02428_),
    .RESET_B(net143),
    .Q(\line_cache[281][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28617_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02429_),
    .RESET_B(net143),
    .Q(\line_cache[281][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28618_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02430_),
    .RESET_B(net143),
    .Q(\line_cache[281][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28619_ (.CLK(clknet_leaf_360_clk_i),
    .D(_02431_),
    .RESET_B(net163),
    .Q(\line_cache[281][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28620_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02432_),
    .RESET_B(net164),
    .Q(\line_cache[281][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28621_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02433_),
    .RESET_B(net164),
    .Q(\line_cache[281][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28622_ (.CLK(clknet_leaf_359_clk_i),
    .D(_02434_),
    .RESET_B(net164),
    .Q(\line_cache[281][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28623_ (.CLK(clknet_leaf_360_clk_i),
    .D(_02435_),
    .RESET_B(net163),
    .Q(\line_cache[282][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28624_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02436_),
    .RESET_B(net141),
    .Q(\line_cache[282][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28625_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02437_),
    .RESET_B(net143),
    .Q(\line_cache[282][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28626_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02438_),
    .RESET_B(net141),
    .Q(\line_cache[282][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28627_ (.CLK(clknet_leaf_359_clk_i),
    .D(_02439_),
    .RESET_B(net163),
    .Q(\line_cache[282][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28628_ (.CLK(clknet_leaf_360_clk_i),
    .D(_02440_),
    .RESET_B(net159),
    .Q(\line_cache[282][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28629_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02441_),
    .RESET_B(net164),
    .Q(\line_cache[282][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28630_ (.CLK(clknet_leaf_359_clk_i),
    .D(_02442_),
    .RESET_B(net163),
    .Q(\line_cache[282][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28631_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02443_),
    .RESET_B(net143),
    .Q(\line_cache[283][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28632_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02444_),
    .RESET_B(net159),
    .Q(\line_cache[283][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28633_ (.CLK(clknet_leaf_363_clk_i),
    .D(_02445_),
    .RESET_B(net143),
    .Q(\line_cache[283][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28634_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02446_),
    .RESET_B(net141),
    .Q(\line_cache[283][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28635_ (.CLK(clknet_leaf_360_clk_i),
    .D(_02447_),
    .RESET_B(net163),
    .Q(\line_cache[283][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28636_ (.CLK(clknet_leaf_359_clk_i),
    .D(_02448_),
    .RESET_B(net163),
    .Q(\line_cache[283][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28637_ (.CLK(clknet_leaf_359_clk_i),
    .D(_02449_),
    .RESET_B(net163),
    .Q(\line_cache[283][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28638_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02450_),
    .RESET_B(net164),
    .Q(\line_cache[283][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28639_ (.CLK(clknet_leaf_361_clk_i),
    .D(_02451_),
    .RESET_B(net163),
    .Q(\line_cache[284][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28640_ (.CLK(clknet_leaf_362_clk_i),
    .D(_02452_),
    .RESET_B(net144),
    .Q(\line_cache[284][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28641_ (.CLK(clknet_leaf_362_clk_i),
    .D(_02453_),
    .RESET_B(net163),
    .Q(\line_cache[284][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28642_ (.CLK(clknet_leaf_362_clk_i),
    .D(_02454_),
    .RESET_B(net144),
    .Q(\line_cache[284][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28643_ (.CLK(clknet_leaf_361_clk_i),
    .D(_02455_),
    .RESET_B(net166),
    .Q(\line_cache[284][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28644_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02456_),
    .RESET_B(net166),
    .Q(\line_cache[284][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28645_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02457_),
    .RESET_B(net165),
    .Q(\line_cache[284][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28646_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02458_),
    .RESET_B(net165),
    .Q(\line_cache[284][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28647_ (.CLK(clknet_leaf_361_clk_i),
    .D(_02459_),
    .RESET_B(net166),
    .Q(\line_cache[285][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28648_ (.CLK(clknet_leaf_30_clk_i),
    .D(_02460_),
    .RESET_B(net175),
    .Q(\line_cache[285][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28649_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02461_),
    .RESET_B(net166),
    .Q(\line_cache[285][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28650_ (.CLK(clknet_leaf_9_clk_i),
    .D(_02462_),
    .RESET_B(net166),
    .Q(\line_cache[285][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28651_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02463_),
    .RESET_B(net166),
    .Q(\line_cache[285][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28652_ (.CLK(clknet_leaf_335_clk_i),
    .D(_02464_),
    .RESET_B(net166),
    .Q(\line_cache[285][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28653_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02465_),
    .RESET_B(net165),
    .Q(\line_cache[285][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28654_ (.CLK(clknet_leaf_334_clk_i),
    .D(_02466_),
    .RESET_B(net176),
    .Q(\line_cache[285][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28655_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02467_),
    .RESET_B(net175),
    .Q(\line_cache[286][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28656_ (.CLK(clknet_leaf_29_clk_i),
    .D(_02468_),
    .RESET_B(net154),
    .Q(\line_cache[286][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28657_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02469_),
    .RESET_B(net154),
    .Q(\line_cache[286][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28658_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02470_),
    .RESET_B(net177),
    .Q(\line_cache[286][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28659_ (.CLK(clknet_leaf_28_clk_i),
    .D(_02471_),
    .RESET_B(net154),
    .Q(\line_cache[286][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28660_ (.CLK(clknet_leaf_31_clk_i),
    .D(_02472_),
    .RESET_B(net177),
    .Q(\line_cache[286][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28661_ (.CLK(clknet_leaf_35_clk_i),
    .D(_02473_),
    .RESET_B(net177),
    .Q(\line_cache[286][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28662_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02474_),
    .RESET_B(net177),
    .Q(\line_cache[286][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28663_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02475_),
    .RESET_B(net176),
    .Q(\line_cache[287][0] ));
 sky130_fd_sc_hd__dfrtp_2 _28664_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02476_),
    .RESET_B(net176),
    .Q(\line_cache[287][1] ));
 sky130_fd_sc_hd__dfrtp_2 _28665_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02477_),
    .RESET_B(net177),
    .Q(\line_cache[287][2] ));
 sky130_fd_sc_hd__dfrtp_2 _28666_ (.CLK(clknet_leaf_333_clk_i),
    .D(_02478_),
    .RESET_B(net177),
    .Q(\line_cache[287][3] ));
 sky130_fd_sc_hd__dfrtp_2 _28667_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02479_),
    .RESET_B(net177),
    .Q(\line_cache[287][4] ));
 sky130_fd_sc_hd__dfrtp_2 _28668_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02480_),
    .RESET_B(net177),
    .Q(\line_cache[287][5] ));
 sky130_fd_sc_hd__dfrtp_2 _28669_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02481_),
    .RESET_B(net177),
    .Q(\line_cache[287][6] ));
 sky130_fd_sc_hd__dfrtp_2 _28670_ (.CLK(clknet_leaf_32_clk_i),
    .D(_02482_),
    .RESET_B(net177),
    .Q(\line_cache[287][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28671_ (.CLK(clknet_leaf_357_clk_i),
    .D(_02483_),
    .RESET_B(net161),
    .Q(\line_cache[288][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28672_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02484_),
    .RESET_B(net161),
    .Q(\line_cache[288][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28673_ (.CLK(clknet_leaf_357_clk_i),
    .D(_02485_),
    .RESET_B(net161),
    .Q(\line_cache[288][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28674_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02486_),
    .RESET_B(net161),
    .Q(\line_cache[288][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28675_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02487_),
    .RESET_B(net167),
    .Q(\line_cache[288][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28676_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02488_),
    .RESET_B(net167),
    .Q(\line_cache[288][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28677_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02489_),
    .RESET_B(net167),
    .Q(\line_cache[288][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28678_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02490_),
    .RESET_B(net167),
    .Q(\line_cache[288][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28679_ (.CLK(clknet_leaf_357_clk_i),
    .D(_02491_),
    .RESET_B(net161),
    .Q(\line_cache[289][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28680_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02492_),
    .RESET_B(net161),
    .Q(\line_cache[289][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28681_ (.CLK(clknet_leaf_351_clk_i),
    .D(_02493_),
    .RESET_B(net162),
    .Q(\line_cache[289][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28682_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02494_),
    .RESET_B(net161),
    .Q(\line_cache[289][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28683_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02495_),
    .RESET_B(net161),
    .Q(\line_cache[289][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28684_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02496_),
    .RESET_B(net167),
    .Q(\line_cache[289][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28685_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02497_),
    .RESET_B(net167),
    .Q(\line_cache[289][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28686_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02498_),
    .RESET_B(net167),
    .Q(\line_cache[289][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28687_ (.CLK(clknet_leaf_351_clk_i),
    .D(_02499_),
    .RESET_B(net162),
    .Q(\line_cache[290][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28688_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02500_),
    .RESET_B(net161),
    .Q(\line_cache[290][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28689_ (.CLK(clknet_leaf_351_clk_i),
    .D(_02501_),
    .RESET_B(net162),
    .Q(\line_cache[290][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28690_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02502_),
    .RESET_B(net161),
    .Q(\line_cache[290][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28691_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02503_),
    .RESET_B(net161),
    .Q(\line_cache[290][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28692_ (.CLK(clknet_leaf_349_clk_i),
    .D(_02504_),
    .RESET_B(net167),
    .Q(\line_cache[290][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28693_ (.CLK(clknet_leaf_349_clk_i),
    .D(_02505_),
    .RESET_B(net167),
    .Q(\line_cache[290][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28694_ (.CLK(clknet_leaf_351_clk_i),
    .D(_02506_),
    .RESET_B(net168),
    .Q(\line_cache[290][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28695_ (.CLK(clknet_leaf_357_clk_i),
    .D(_02507_),
    .RESET_B(net162),
    .Q(\line_cache[291][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28696_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02508_),
    .RESET_B(net161),
    .Q(\line_cache[291][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28697_ (.CLK(clknet_leaf_351_clk_i),
    .D(_02509_),
    .RESET_B(net162),
    .Q(\line_cache[291][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28698_ (.CLK(clknet_leaf_352_clk_i),
    .D(_02510_),
    .RESET_B(net161),
    .Q(\line_cache[291][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28699_ (.CLK(clknet_leaf_349_clk_i),
    .D(_02511_),
    .RESET_B(net167),
    .Q(\line_cache[291][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28700_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02512_),
    .RESET_B(net167),
    .Q(\line_cache[291][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28701_ (.CLK(clknet_leaf_349_clk_i),
    .D(_02513_),
    .RESET_B(net167),
    .Q(\line_cache[291][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28702_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02514_),
    .RESET_B(net168),
    .Q(\line_cache[291][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28703_ (.CLK(clknet_leaf_356_clk_i),
    .D(_02515_),
    .RESET_B(net159),
    .Q(\line_cache[292][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28704_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02516_),
    .RESET_B(net159),
    .Q(\line_cache[292][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28705_ (.CLK(clknet_leaf_356_clk_i),
    .D(_02517_),
    .RESET_B(net159),
    .Q(\line_cache[292][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28706_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02518_),
    .RESET_B(net159),
    .Q(\line_cache[292][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28707_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02519_),
    .RESET_B(net161),
    .Q(\line_cache[292][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28708_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02520_),
    .RESET_B(net161),
    .Q(\line_cache[292][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28709_ (.CLK(clknet_leaf_357_clk_i),
    .D(_02521_),
    .RESET_B(net162),
    .Q(\line_cache[292][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28710_ (.CLK(clknet_leaf_357_clk_i),
    .D(_02522_),
    .RESET_B(net162),
    .Q(\line_cache[292][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28711_ (.CLK(clknet_leaf_356_clk_i),
    .D(_02523_),
    .RESET_B(net160),
    .Q(\line_cache[293][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28712_ (.CLK(clknet_leaf_354_clk_i),
    .D(_02524_),
    .RESET_B(net159),
    .Q(\line_cache[293][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28713_ (.CLK(clknet_leaf_356_clk_i),
    .D(_02525_),
    .RESET_B(net160),
    .Q(\line_cache[293][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28714_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02526_),
    .RESET_B(net159),
    .Q(\line_cache[293][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28715_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02527_),
    .RESET_B(net161),
    .Q(\line_cache[293][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28716_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02528_),
    .RESET_B(net159),
    .Q(\line_cache[293][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28717_ (.CLK(clknet_leaf_355_clk_i),
    .D(_02529_),
    .RESET_B(net160),
    .Q(\line_cache[293][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28718_ (.CLK(clknet_leaf_356_clk_i),
    .D(_02530_),
    .RESET_B(net160),
    .Q(\line_cache[293][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28719_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02531_),
    .RESET_B(net141),
    .Q(\line_cache[294][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28720_ (.CLK(clknet_leaf_366_clk_i),
    .D(_02532_),
    .RESET_B(net159),
    .Q(\line_cache[294][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28721_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02533_),
    .RESET_B(net145),
    .Q(\line_cache[294][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28722_ (.CLK(clknet_leaf_354_clk_i),
    .D(_02534_),
    .RESET_B(net159),
    .Q(\line_cache[294][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28723_ (.CLK(clknet_leaf_366_clk_i),
    .D(_02535_),
    .RESET_B(net159),
    .Q(\line_cache[294][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28724_ (.CLK(clknet_leaf_354_clk_i),
    .D(_02536_),
    .RESET_B(net159),
    .Q(\line_cache[294][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28725_ (.CLK(clknet_leaf_355_clk_i),
    .D(_02537_),
    .RESET_B(net160),
    .Q(\line_cache[294][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28726_ (.CLK(clknet_leaf_355_clk_i),
    .D(_02538_),
    .RESET_B(net160),
    .Q(\line_cache[294][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28727_ (.CLK(clknet_leaf_356_clk_i),
    .D(_02539_),
    .RESET_B(net160),
    .Q(\line_cache[295][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28728_ (.CLK(clknet_leaf_354_clk_i),
    .D(_02540_),
    .RESET_B(net159),
    .Q(\line_cache[295][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28729_ (.CLK(clknet_leaf_365_clk_i),
    .D(_02541_),
    .RESET_B(net145),
    .Q(\line_cache[295][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28730_ (.CLK(clknet_leaf_353_clk_i),
    .D(_02542_),
    .RESET_B(net159),
    .Q(\line_cache[295][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28731_ (.CLK(clknet_leaf_366_clk_i),
    .D(_02543_),
    .RESET_B(net141),
    .Q(\line_cache[295][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28732_ (.CLK(clknet_leaf_354_clk_i),
    .D(_02544_),
    .RESET_B(net159),
    .Q(\line_cache[295][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28733_ (.CLK(clknet_leaf_355_clk_i),
    .D(_02545_),
    .RESET_B(net160),
    .Q(\line_cache[295][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28734_ (.CLK(clknet_leaf_355_clk_i),
    .D(_02546_),
    .RESET_B(net160),
    .Q(\line_cache[295][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28735_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02547_),
    .RESET_B(net164),
    .Q(\line_cache[296][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28736_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02548_),
    .RESET_B(net164),
    .Q(\line_cache[296][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28737_ (.CLK(clknet_leaf_338_clk_i),
    .D(_02549_),
    .RESET_B(net172),
    .Q(\line_cache[296][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28738_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02550_),
    .RESET_B(net164),
    .Q(\line_cache[296][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28739_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02551_),
    .RESET_B(net171),
    .Q(\line_cache[296][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28740_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02552_),
    .RESET_B(net171),
    .Q(\line_cache[296][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28741_ (.CLK(clknet_leaf_339_clk_i),
    .D(_02553_),
    .RESET_B(net172),
    .Q(\line_cache[296][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28742_ (.CLK(clknet_leaf_338_clk_i),
    .D(_02554_),
    .RESET_B(net172),
    .Q(\line_cache[296][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28743_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02555_),
    .RESET_B(net164),
    .Q(\line_cache[297][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28744_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02556_),
    .RESET_B(net164),
    .Q(\line_cache[297][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28745_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02557_),
    .RESET_B(net165),
    .Q(\line_cache[297][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28746_ (.CLK(clknet_leaf_358_clk_i),
    .D(_02558_),
    .RESET_B(net162),
    .Q(\line_cache[297][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28747_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02559_),
    .RESET_B(net171),
    .Q(\line_cache[297][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28748_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02560_),
    .RESET_B(net172),
    .Q(\line_cache[297][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28749_ (.CLK(clknet_leaf_338_clk_i),
    .D(_02561_),
    .RESET_B(net172),
    .Q(\line_cache[297][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28750_ (.CLK(clknet_leaf_338_clk_i),
    .D(_02562_),
    .RESET_B(net172),
    .Q(\line_cache[297][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28751_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02563_),
    .RESET_B(net171),
    .Q(\line_cache[298][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28752_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02564_),
    .RESET_B(net171),
    .Q(\line_cache[298][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28753_ (.CLK(clknet_leaf_336_clk_i),
    .D(_02565_),
    .RESET_B(net165),
    .Q(\line_cache[298][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28754_ (.CLK(clknet_leaf_351_clk_i),
    .D(_02566_),
    .RESET_B(net168),
    .Q(\line_cache[298][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28755_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02567_),
    .RESET_B(net168),
    .Q(\line_cache[298][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28756_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02568_),
    .RESET_B(net171),
    .Q(\line_cache[298][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28757_ (.CLK(clknet_leaf_338_clk_i),
    .D(_02569_),
    .RESET_B(net171),
    .Q(\line_cache[298][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28758_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02570_),
    .RESET_B(net171),
    .Q(\line_cache[298][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28759_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02571_),
    .RESET_B(net171),
    .Q(\line_cache[299][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28760_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02572_),
    .RESET_B(net171),
    .Q(\line_cache[299][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28761_ (.CLK(clknet_leaf_338_clk_i),
    .D(_02573_),
    .RESET_B(net172),
    .Q(\line_cache[299][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28762_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02574_),
    .RESET_B(net168),
    .Q(\line_cache[299][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28763_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02575_),
    .RESET_B(net168),
    .Q(\line_cache[299][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28764_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02576_),
    .RESET_B(net172),
    .Q(\line_cache[299][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28765_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02577_),
    .RESET_B(net172),
    .Q(\line_cache[299][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28766_ (.CLK(clknet_leaf_337_clk_i),
    .D(_02578_),
    .RESET_B(net171),
    .Q(\line_cache[299][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28767_ (.CLK(clknet_leaf_342_clk_i),
    .D(_02579_),
    .RESET_B(net248),
    .Q(\line_cache[300][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28768_ (.CLK(clknet_leaf_342_clk_i),
    .D(_02580_),
    .RESET_B(net172),
    .Q(\line_cache[300][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28769_ (.CLK(clknet_leaf_342_clk_i),
    .D(_02581_),
    .RESET_B(net172),
    .Q(\line_cache[300][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28770_ (.CLK(clknet_leaf_342_clk_i),
    .D(_02582_),
    .RESET_B(net172),
    .Q(\line_cache[300][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28771_ (.CLK(clknet_leaf_342_clk_i),
    .D(_02583_),
    .RESET_B(net172),
    .Q(\line_cache[300][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28772_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02584_),
    .RESET_B(net248),
    .Q(\line_cache[300][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28773_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02585_),
    .RESET_B(net248),
    .Q(\line_cache[300][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28774_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02586_),
    .RESET_B(net248),
    .Q(\line_cache[300][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28775_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02587_),
    .RESET_B(net248),
    .Q(\line_cache[301][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28776_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02588_),
    .RESET_B(net173),
    .Q(\line_cache[301][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28777_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02589_),
    .RESET_B(net173),
    .Q(\line_cache[301][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28778_ (.CLK(clknet_leaf_341_clk_i),
    .D(_02590_),
    .RESET_B(net173),
    .Q(\line_cache[301][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28779_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02591_),
    .RESET_B(net173),
    .Q(\line_cache[301][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28780_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02592_),
    .RESET_B(net248),
    .Q(\line_cache[301][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28781_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02593_),
    .RESET_B(net250),
    .Q(\line_cache[301][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28782_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02594_),
    .RESET_B(net250),
    .Q(\line_cache[301][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28783_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02595_),
    .RESET_B(net258),
    .Q(\line_cache[302][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28784_ (.CLK(clknet_leaf_331_clk_i),
    .D(_02596_),
    .RESET_B(net182),
    .Q(\line_cache[302][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28785_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02597_),
    .RESET_B(net173),
    .Q(\line_cache[302][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28786_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02598_),
    .RESET_B(net182),
    .Q(\line_cache[302][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28787_ (.CLK(clknet_leaf_340_clk_i),
    .D(_02599_),
    .RESET_B(net173),
    .Q(\line_cache[302][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28788_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02600_),
    .RESET_B(net250),
    .Q(\line_cache[302][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28789_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02601_),
    .RESET_B(net250),
    .Q(\line_cache[302][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28790_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02602_),
    .RESET_B(net250),
    .Q(\line_cache[302][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28791_ (.CLK(clknet_leaf_321_clk_i),
    .D(_02603_),
    .RESET_B(net258),
    .Q(\line_cache[303][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28792_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02604_),
    .RESET_B(net258),
    .Q(\line_cache[303][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28793_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02605_),
    .RESET_B(net250),
    .Q(\line_cache[303][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28794_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02606_),
    .RESET_B(net258),
    .Q(\line_cache[303][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28795_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02607_),
    .RESET_B(net258),
    .Q(\line_cache[303][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28796_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02608_),
    .RESET_B(net262),
    .Q(\line_cache[303][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28797_ (.CLK(clknet_leaf_320_clk_i),
    .D(_02609_),
    .RESET_B(net258),
    .Q(\line_cache[303][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28798_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02610_),
    .RESET_B(net250),
    .Q(\line_cache[303][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28799_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02611_),
    .RESET_B(net244),
    .Q(\line_cache[304][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28800_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02612_),
    .RESET_B(net244),
    .Q(\line_cache[304][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28801_ (.CLK(clknet_leaf_345_clk_i),
    .D(_02613_),
    .RESET_B(net169),
    .Q(\line_cache[304][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28802_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02614_),
    .RESET_B(net246),
    .Q(\line_cache[304][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28803_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02615_),
    .RESET_B(net251),
    .Q(\line_cache[304][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28804_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02616_),
    .RESET_B(net251),
    .Q(\line_cache[304][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28805_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02617_),
    .RESET_B(net246),
    .Q(\line_cache[304][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28806_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02618_),
    .RESET_B(net244),
    .Q(\line_cache[304][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28807_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02619_),
    .RESET_B(net244),
    .Q(\line_cache[305][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28808_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02620_),
    .RESET_B(net244),
    .Q(\line_cache[305][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28809_ (.CLK(clknet_leaf_303_clk_i),
    .D(_02621_),
    .RESET_B(net244),
    .Q(\line_cache[305][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28810_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02622_),
    .RESET_B(net246),
    .Q(\line_cache[305][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28811_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02623_),
    .RESET_B(net246),
    .Q(\line_cache[305][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28812_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02624_),
    .RESET_B(net246),
    .Q(\line_cache[305][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28813_ (.CLK(clknet_leaf_297_clk_i),
    .D(_02625_),
    .RESET_B(net246),
    .Q(\line_cache[305][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28814_ (.CLK(clknet_leaf_303_clk_i),
    .D(_02626_),
    .RESET_B(net244),
    .Q(\line_cache[305][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28815_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02627_),
    .RESET_B(net244),
    .Q(\line_cache[306][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28816_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02628_),
    .RESET_B(net244),
    .Q(\line_cache[306][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28817_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02629_),
    .RESET_B(net244),
    .Q(\line_cache[306][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28818_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02630_),
    .RESET_B(net246),
    .Q(\line_cache[306][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28819_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02631_),
    .RESET_B(net251),
    .Q(\line_cache[306][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28820_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02632_),
    .RESET_B(net251),
    .Q(\line_cache[306][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28821_ (.CLK(clknet_leaf_296_clk_i),
    .D(_02633_),
    .RESET_B(net246),
    .Q(\line_cache[306][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28822_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02634_),
    .RESET_B(net244),
    .Q(\line_cache[306][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28823_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02635_),
    .RESET_B(net244),
    .Q(\line_cache[307][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28824_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02636_),
    .RESET_B(net244),
    .Q(\line_cache[307][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28825_ (.CLK(clknet_leaf_302_clk_i),
    .D(_02637_),
    .RESET_B(net244),
    .Q(\line_cache[307][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28826_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02638_),
    .RESET_B(net246),
    .Q(\line_cache[307][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28827_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02639_),
    .RESET_B(net246),
    .Q(\line_cache[307][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28828_ (.CLK(clknet_leaf_300_clk_i),
    .D(_02640_),
    .RESET_B(net246),
    .Q(\line_cache[307][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28829_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02641_),
    .RESET_B(net246),
    .Q(\line_cache[307][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28830_ (.CLK(clknet_leaf_301_clk_i),
    .D(_02642_),
    .RESET_B(net244),
    .Q(\line_cache[307][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28831_ (.CLK(clknet_leaf_345_clk_i),
    .D(_02643_),
    .RESET_B(net169),
    .Q(\line_cache[308][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28832_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02644_),
    .RESET_B(net169),
    .Q(\line_cache[308][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28833_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02645_),
    .RESET_B(net173),
    .Q(\line_cache[308][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28834_ (.CLK(clknet_leaf_347_clk_i),
    .D(_02646_),
    .RESET_B(net169),
    .Q(\line_cache[308][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28835_ (.CLK(clknet_leaf_347_clk_i),
    .D(_02647_),
    .RESET_B(net169),
    .Q(\line_cache[308][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28836_ (.CLK(clknet_leaf_347_clk_i),
    .D(_02648_),
    .RESET_B(net169),
    .Q(\line_cache[308][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28837_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02649_),
    .RESET_B(net169),
    .Q(\line_cache[308][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28838_ (.CLK(clknet_leaf_345_clk_i),
    .D(_02650_),
    .RESET_B(net169),
    .Q(\line_cache[308][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28839_ (.CLK(clknet_leaf_345_clk_i),
    .D(_02651_),
    .RESET_B(net170),
    .Q(\line_cache[309][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28840_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02652_),
    .RESET_B(net169),
    .Q(\line_cache[309][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28841_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02653_),
    .RESET_B(net170),
    .Q(\line_cache[309][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28842_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02654_),
    .RESET_B(net167),
    .Q(\line_cache[309][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28843_ (.CLK(clknet_leaf_347_clk_i),
    .D(_02655_),
    .RESET_B(net169),
    .Q(\line_cache[309][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28844_ (.CLK(clknet_leaf_347_clk_i),
    .D(_02656_),
    .RESET_B(net169),
    .Q(\line_cache[309][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28845_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02657_),
    .RESET_B(net169),
    .Q(\line_cache[309][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28846_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02658_),
    .RESET_B(net170),
    .Q(\line_cache[309][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28847_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02659_),
    .RESET_B(net168),
    .Q(\line_cache[310][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28848_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02660_),
    .RESET_B(net168),
    .Q(\line_cache[310][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28849_ (.CLK(clknet_leaf_345_clk_i),
    .D(_02661_),
    .RESET_B(net170),
    .Q(\line_cache[310][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28850_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02662_),
    .RESET_B(net167),
    .Q(\line_cache[310][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28851_ (.CLK(clknet_leaf_347_clk_i),
    .D(_02663_),
    .RESET_B(net169),
    .Q(\line_cache[310][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28852_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02664_),
    .RESET_B(net169),
    .Q(\line_cache[310][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28853_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02665_),
    .RESET_B(net170),
    .Q(\line_cache[310][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28854_ (.CLK(clknet_leaf_350_clk_i),
    .D(_02666_),
    .RESET_B(net168),
    .Q(\line_cache[310][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28855_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02667_),
    .RESET_B(net168),
    .Q(\line_cache[311][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28856_ (.CLK(clknet_leaf_349_clk_i),
    .D(_02668_),
    .RESET_B(net167),
    .Q(\line_cache[311][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28857_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02669_),
    .RESET_B(net170),
    .Q(\line_cache[311][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28858_ (.CLK(clknet_leaf_348_clk_i),
    .D(_02670_),
    .RESET_B(net167),
    .Q(\line_cache[311][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28859_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02671_),
    .RESET_B(net169),
    .Q(\line_cache[311][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28860_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02672_),
    .RESET_B(net169),
    .Q(\line_cache[311][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28861_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02673_),
    .RESET_B(net170),
    .Q(\line_cache[311][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28862_ (.CLK(clknet_leaf_344_clk_i),
    .D(_02674_),
    .RESET_B(net168),
    .Q(\line_cache[311][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28863_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02675_),
    .RESET_B(net173),
    .Q(\line_cache[312][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28864_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02676_),
    .RESET_B(net170),
    .Q(\line_cache[312][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28865_ (.CLK(clknet_leaf_345_clk_i),
    .D(_02677_),
    .RESET_B(net170),
    .Q(\line_cache[312][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28866_ (.CLK(clknet_leaf_299_clk_i),
    .D(_02678_),
    .RESET_B(net246),
    .Q(\line_cache[312][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28867_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02679_),
    .RESET_B(net246),
    .Q(\line_cache[312][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28868_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02680_),
    .RESET_B(net246),
    .Q(\line_cache[312][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28869_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02681_),
    .RESET_B(net249),
    .Q(\line_cache[312][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28870_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02682_),
    .RESET_B(net248),
    .Q(\line_cache[312][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28871_ (.CLK(clknet_leaf_343_clk_i),
    .D(_02683_),
    .RESET_B(net244),
    .Q(\line_cache[313][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28872_ (.CLK(clknet_leaf_303_clk_i),
    .D(_02684_),
    .RESET_B(net245),
    .Q(\line_cache[313][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28873_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02685_),
    .RESET_B(net245),
    .Q(\line_cache[313][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28874_ (.CLK(clknet_leaf_303_clk_i),
    .D(_02686_),
    .RESET_B(net245),
    .Q(\line_cache[313][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28875_ (.CLK(clknet_leaf_298_clk_i),
    .D(_02687_),
    .RESET_B(net246),
    .Q(\line_cache[313][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28876_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02688_),
    .RESET_B(net247),
    .Q(\line_cache[313][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28877_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02689_),
    .RESET_B(net249),
    .Q(\line_cache[313][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28878_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02690_),
    .RESET_B(net248),
    .Q(\line_cache[313][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28879_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02691_),
    .RESET_B(net248),
    .Q(\line_cache[314][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28880_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02692_),
    .RESET_B(net245),
    .Q(\line_cache[314][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28881_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02693_),
    .RESET_B(net245),
    .Q(\line_cache[314][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28882_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02694_),
    .RESET_B(net247),
    .Q(\line_cache[314][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28883_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02695_),
    .RESET_B(net247),
    .Q(\line_cache[314][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28884_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02696_),
    .RESET_B(net247),
    .Q(\line_cache[314][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28885_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02697_),
    .RESET_B(net249),
    .Q(\line_cache[314][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28886_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02698_),
    .RESET_B(net248),
    .Q(\line_cache[314][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28887_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02699_),
    .RESET_B(net248),
    .Q(\line_cache[315][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28888_ (.CLK(clknet_leaf_346_clk_i),
    .D(_02700_),
    .RESET_B(net245),
    .Q(\line_cache[315][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28889_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02701_),
    .RESET_B(net245),
    .Q(\line_cache[315][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28890_ (.CLK(clknet_leaf_304_clk_i),
    .D(_02702_),
    .RESET_B(net245),
    .Q(\line_cache[315][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28891_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02703_),
    .RESET_B(net247),
    .Q(\line_cache[315][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28892_ (.CLK(clknet_leaf_305_clk_i),
    .D(_02704_),
    .RESET_B(net247),
    .Q(\line_cache[315][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28893_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02705_),
    .RESET_B(net249),
    .Q(\line_cache[315][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28894_ (.CLK(clknet_leaf_307_clk_i),
    .D(_02706_),
    .RESET_B(net248),
    .Q(\line_cache[315][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28895_ (.CLK(clknet_leaf_309_clk_i),
    .D(_02707_),
    .RESET_B(net249),
    .Q(\line_cache[316][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28896_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02708_),
    .RESET_B(net248),
    .Q(\line_cache[316][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28897_ (.CLK(clknet_leaf_306_clk_i),
    .D(_02709_),
    .RESET_B(net249),
    .Q(\line_cache[316][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28898_ (.CLK(clknet_leaf_308_clk_i),
    .D(_02710_),
    .RESET_B(net248),
    .Q(\line_cache[316][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28899_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02711_),
    .RESET_B(net249),
    .Q(\line_cache[316][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28900_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02712_),
    .RESET_B(net249),
    .Q(\line_cache[316][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28901_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02713_),
    .RESET_B(net249),
    .Q(\line_cache[316][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28902_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02714_),
    .RESET_B(net249),
    .Q(\line_cache[316][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28903_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02715_),
    .RESET_B(net249),
    .Q(\line_cache[317][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28904_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02716_),
    .RESET_B(net249),
    .Q(\line_cache[317][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28905_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02717_),
    .RESET_B(net249),
    .Q(\line_cache[317][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28906_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02718_),
    .RESET_B(net250),
    .Q(\line_cache[317][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28907_ (.CLK(clknet_leaf_312_clk_i),
    .D(_02719_),
    .RESET_B(net249),
    .Q(\line_cache[317][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28908_ (.CLK(clknet_leaf_313_clk_i),
    .D(_02720_),
    .RESET_B(net249),
    .Q(\line_cache[317][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28909_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02721_),
    .RESET_B(net250),
    .Q(\line_cache[317][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28910_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02722_),
    .RESET_B(net250),
    .Q(\line_cache[317][7] ));
 sky130_fd_sc_hd__dfrtp_1 _28911_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02723_),
    .RESET_B(net250),
    .Q(\line_cache[318][0] ));
 sky130_fd_sc_hd__dfrtp_1 _28912_ (.CLK(clknet_leaf_319_clk_i),
    .D(_02724_),
    .RESET_B(net262),
    .Q(\line_cache[318][1] ));
 sky130_fd_sc_hd__dfrtp_1 _28913_ (.CLK(clknet_leaf_310_clk_i),
    .D(_02725_),
    .RESET_B(net250),
    .Q(\line_cache[318][2] ));
 sky130_fd_sc_hd__dfrtp_1 _28914_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02726_),
    .RESET_B(net257),
    .Q(\line_cache[318][3] ));
 sky130_fd_sc_hd__dfrtp_1 _28915_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02727_),
    .RESET_B(net250),
    .Q(\line_cache[318][4] ));
 sky130_fd_sc_hd__dfrtp_1 _28916_ (.CLK(clknet_leaf_311_clk_i),
    .D(_02728_),
    .RESET_B(net250),
    .Q(\line_cache[318][5] ));
 sky130_fd_sc_hd__dfrtp_1 _28917_ (.CLK(clknet_leaf_319_clk_i),
    .D(_02729_),
    .RESET_B(net263),
    .Q(\line_cache[318][6] ));
 sky130_fd_sc_hd__dfrtp_1 _28918_ (.CLK(clknet_leaf_319_clk_i),
    .D(_02730_),
    .RESET_B(net263),
    .Q(\line_cache[318][7] ));
 sky130_fd_sc_hd__dfrtp_2 _28919_ (.CLK(clknet_leaf_275_clk_i),
    .D(_02731_),
    .RESET_B(net279),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _28920_ (.CLK(clknet_leaf_366_clk_i),
    .D(_02732_),
    .RESET_B(net141),
    .Q(net123));
 sky130_fd_sc_hd__buf_1 _28957_ (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_0_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_1_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_2_0_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_3_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_10__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_11__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_12__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_13__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_14__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_15__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_16__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_17__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_18__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_19__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_20__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_21__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_22__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk_i (.A(clknet_2_2_0_clk_i),
    .X(clknet_5_23__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_24__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_25__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_26__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_27__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_28__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_29__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_30__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk_i (.A(clknet_2_3_0_clk_i),
    .X(clknet_5_31__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_3__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_4__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_5__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_6__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk_i (.A(clknet_2_0_0_clk_i),
    .X(clknet_5_7__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_8__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk_i (.A(clknet_2_1_0_clk_i),
    .X(clknet_5_9__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_100_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_101_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_102_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_103_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_104_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_105_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_106_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_107_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_108_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_109_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_110_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_111_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_112_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_113_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_114_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_115_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_116_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_117_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_118_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_119_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_120_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_121_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_122_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk_i (.A(clknet_5_15__leaf_clk_i),
    .X(clknet_leaf_123_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_124_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_125_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_126_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk_i (.A(clknet_5_14__leaf_clk_i),
    .X(clknet_leaf_127_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_128_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_129_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_130_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_131_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_132_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_133_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_134_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_135_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_136_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_137_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_138_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_139_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_140_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_141_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_142_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_143_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_144_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_145_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_146_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_147_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_148_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_149_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_150_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_151_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_152_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_153_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_154_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_155_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_156_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_157_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_158_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_159_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_160_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_161_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_162_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_163_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_164_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk_i (.A(clknet_5_26__leaf_clk_i),
    .X(clknet_leaf_165_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_166_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_167_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_168_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_169_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_170_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_171_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_172_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_173_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_174_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_175_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_176_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_177_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_178_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_179_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_180_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_181_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_182_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_183_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_184_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_185_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_186_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_187_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_188_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_189_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_190_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk_i (.A(clknet_5_27__leaf_clk_i),
    .X(clknet_leaf_191_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk_i (.A(clknet_5_30__leaf_clk_i),
    .X(clknet_leaf_192_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_193_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_194_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_195_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_196_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk_i (.A(clknet_5_31__leaf_clk_i),
    .X(clknet_leaf_197_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_198_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_199_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_200_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_201_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_202_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_203_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_204_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_205_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_206_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_207_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_208_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_209_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_210_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_211_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_212_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_213_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_214_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_215_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_216_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_217_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_218_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_219_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_220_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_221_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_222_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_223_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_224_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_225_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_226_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_227_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_228_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk_i (.A(clknet_5_24__leaf_clk_i),
    .X(clknet_leaf_229_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_230_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_231_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk_i (.A(clknet_5_25__leaf_clk_i),
    .X(clknet_leaf_232_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_233_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_234_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_235_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_236_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_237_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_238_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_239_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_240_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_241_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_242_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_243_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_244_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_245_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_246_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_247_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk_i (.A(clknet_5_28__leaf_clk_i),
    .X(clknet_leaf_248_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_249_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_250_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_251_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_252_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk_i (.A(clknet_5_29__leaf_clk_i),
    .X(clknet_leaf_253_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_254_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_255_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_256_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_257_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_258_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_259_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_260_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk_i (.A(clknet_5_23__leaf_clk_i),
    .X(clknet_leaf_261_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_262_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk_i (.A(clknet_5_22__leaf_clk_i),
    .X(clknet_leaf_263_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_264_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_265_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_266_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_267_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_268_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_269_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_270_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_271_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_272_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_273_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_274_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_275_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_276_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk_i (.A(clknet_5_21__leaf_clk_i),
    .X(clknet_leaf_277_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_278_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_279_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_280_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_281_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_282_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_283_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_284_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_285_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_286_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_287_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_288_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_289_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_290_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_291_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_clk_i (.A(clknet_5_20__leaf_clk_i),
    .X(clknet_leaf_292_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_293_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_294_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_295_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_296_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_297_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_298_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_299_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_300_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_301_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_302_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_303_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_304_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_305_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_306_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_306_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_307_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_307_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_308_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_309_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_310_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_311_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_312_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_313_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_clk_i (.A(clknet_5_17__leaf_clk_i),
    .X(clknet_leaf_314_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_315_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_316_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_317_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_318_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_clk_i (.A(clknet_5_19__leaf_clk_i),
    .X(clknet_leaf_319_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_320_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_321_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_322_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_323_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_323_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_324_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_324_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_325_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_325_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_326_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_326_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_327_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_327_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_328_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_328_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_329_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_329_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_330_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_330_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_331_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_331_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_332_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_332_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_333_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_333_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_334_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_334_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_335_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_335_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_336_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_336_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_337_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_337_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_338_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_338_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_339_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_339_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_340_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_340_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_341_clk_i (.A(clknet_5_18__leaf_clk_i),
    .X(clknet_leaf_341_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_342_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_342_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_343_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_343_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_344_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_344_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_345_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_345_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_346_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_346_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_347_clk_i (.A(clknet_5_16__leaf_clk_i),
    .X(clknet_leaf_347_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_348_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_348_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_349_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_349_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_350_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_350_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_351_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_351_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_352_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_352_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_353_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_353_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_354_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_354_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_355_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_355_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_356_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_356_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_357_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_357_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_358_clk_i (.A(clknet_5_5__leaf_clk_i),
    .X(clknet_leaf_358_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_359_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_359_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_360_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_360_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_361_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_361_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_362_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_362_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_363_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_363_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_364_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_364_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_365_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_365_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_366_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_366_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_367_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_367_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_368_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_368_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_370_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_370_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_371_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_371_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_39_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_42_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i (.A(clknet_5_13__leaf_clk_i),
    .X(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_45_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_i (.A(clknet_5_7__leaf_clk_i),
    .X(clknet_leaf_46_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_i (.A(clknet_5_6__leaf_clk_i),
    .X(clknet_leaf_47_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_48_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_49_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_5_0__leaf_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_50_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_51_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_52_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_i (.A(clknet_5_12__leaf_clk_i),
    .X(clknet_leaf_53_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_54_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_55_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_56_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_57_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_58_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_59_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_60_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_i (.A(clknet_5_3__leaf_clk_i),
    .X(clknet_leaf_61_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_62_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_63_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_64_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_65_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_66_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_i (.A(clknet_5_2__leaf_clk_i),
    .X(clknet_leaf_67_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_68_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_69_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_70_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_71_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_72_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_73_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_74_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_75_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_76_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_i (.A(clknet_5_8__leaf_clk_i),
    .X(clknet_leaf_77_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_78_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_79_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_5_1__leaf_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_i (.A(clknet_5_9__leaf_clk_i),
    .X(clknet_leaf_80_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_81_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_82_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_83_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_84_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_85_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_86_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_87_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_88_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_89_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_90_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_91_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_92_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_93_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_i (.A(clknet_5_10__leaf_clk_i),
    .X(clknet_leaf_94_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_95_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_96_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_97_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_98_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_i (.A(clknet_5_11__leaf_clk_i),
    .X(clknet_leaf_99_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_5_4__leaf_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout137 (.A(net146),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net146),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net146),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 fanout140 (.A(net145),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_8 fanout141 (.A(net145),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_8 fanout142 (.A(net145),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net145),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net243),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_8 fanout147 (.A(net158),
    .X(net147));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net158),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_8 fanout149 (.A(net158),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(net158),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_8 fanout151 (.A(net158),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net158),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_8 fanout153 (.A(net158),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net158),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_8 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net243),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_8 fanout159 (.A(net174),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net174),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_8 fanout161 (.A(net174),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net174),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(net166),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__buf_2 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net174),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net174),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net174),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net174),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(net174),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_8 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net243),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(net177),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net243),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_8 fanout178 (.A(net180),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net243),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(net185),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net185),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net243),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(net214),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net214),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net214),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net214),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout190 (.A(net193),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net214),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(net197),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(net197),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net214),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net201),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(net201),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net214),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(net205),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net214),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_8 fanout207 (.A(net214),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(net210),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(net214),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net213),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_8 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_8 fanout214 (.A(net243),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 fanout215 (.A(net217),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_8 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net243),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(net221),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_8 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net243),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_8 fanout222 (.A(net224),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net243),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(net227),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_8 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net243),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_8 fanout228 (.A(net230),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net242),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 fanout231 (.A(net242),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net242),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 fanout233 (.A(net242),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net242),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_8 fanout235 (.A(net242),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(net242),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_8 fanout238 (.A(net241),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net241),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_8 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_8 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_16 fanout243 (.A(net83),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_8 fanout244 (.A(net247),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 fanout245 (.A(net247),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_8 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 fanout247 (.A(net300),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_8 fanout248 (.A(net250),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_8 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_8 fanout250 (.A(net300),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_8 fanout251 (.A(net254),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net254),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 fanout254 (.A(net300),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_8 fanout255 (.A(net257),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(net300),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_8 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 fanout259 (.A(net262),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_8 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(net300),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_8 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 fanout264 (.A(net268),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_8 fanout265 (.A(net267),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_8 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_8 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout268 (.A(net300),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_8 fanout269 (.A(net283),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net283),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_8 fanout271 (.A(net283),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net283),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_8 fanout273 (.A(net276),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_8 fanout274 (.A(net276),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net283),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_8 fanout277 (.A(net279),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_8 fanout279 (.A(net283),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_8 fanout280 (.A(net283),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_8 fanout281 (.A(net283),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_8 fanout283 (.A(net300),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_8 fanout284 (.A(net287),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net300),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_8 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 fanout289 (.A(net291),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net300),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_8 fanout292 (.A(net295),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_8 fanout293 (.A(net295),
    .X(net293));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 fanout295 (.A(net300),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_8 fanout296 (.A(net299),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_8 fanout297 (.A(net299),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_6 fanout300 (.A(net83),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 fanout301 (.A(net303),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_8 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_8 fanout303 (.A(net315),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_8 fanout304 (.A(net315),
    .X(net304));
 sky130_fd_sc_hd__buf_4 fanout305 (.A(net315),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_8 fanout306 (.A(net315),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_8 fanout307 (.A(net315),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(net315),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_8 fanout309 (.A(net315),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net315),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_8 fanout311 (.A(net314),
    .X(net311));
 sky130_fd_sc_hd__buf_4 fanout312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_8 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_8 fanout315 (.A(net353),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_8 fanout316 (.A(net318),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_8 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(net353),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_8 fanout319 (.A(net321),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_8 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_8 fanout321 (.A(net353),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_8 fanout322 (.A(net325),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(net325),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_8 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net353),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_8 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_8 fanout327 (.A(net353),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_8 fanout328 (.A(net331),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_8 fanout329 (.A(net331),
    .X(net329));
 sky130_fd_sc_hd__buf_4 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 fanout331 (.A(net342),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 fanout332 (.A(net334),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_8 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(net342),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_8 fanout335 (.A(net338),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_4 fanout336 (.A(net338),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_8 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 fanout338 (.A(net342),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_8 fanout339 (.A(net342),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net342),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_8 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(net353),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_8 fanout343 (.A(net345),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_8 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_8 fanout345 (.A(net352),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_8 fanout346 (.A(net352),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_8 fanout347 (.A(net352),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_8 fanout348 (.A(net350),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_8 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_8 fanout350 (.A(net352),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_8 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_4 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__buf_4 fanout353 (.A(net83),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\line_cache[105][6] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_02945_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_07925_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_07837_),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\line_cache[102][0] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_04816_),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\line_cache[153][7] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_05836_),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\line_cache[238][1] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_07378_),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\line_cache[206][6] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_06810_),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\line_cache[165][1] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\line_cache[257][5] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_06039_),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\line_cache[91][6] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_04625_),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\line_cache[135][0] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_05456_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\line_cache[265][1] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_07873_),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\line_cache[170][6] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_06146_),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\line_cache[141][1] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_07738_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_05592_),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\line_cache[150][4] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_05774_),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\line_cache[189][0] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_06473_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\line_cache[91][0] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_04613_),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\line_cache[94][6] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_04682_),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\line_cache[238][5] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\line_cache[241][1] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_07387_),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\line_cache[270][0] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_07967_),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\line_cache[70][0] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_04225_),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\line_cache[151][4] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_05791_),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\line_cache[90][6] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_04609_),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\line_cache[141][2] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_07428_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_05596_),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\line_cache[263][3] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_07844_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\line_cache[222][5] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_07098_),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\line_cache[110][6] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_04976_),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\line_cache[90][1] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_04597_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\line_cache[127][5] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\line_cache[105][7] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_05313_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\line_cache[154][5] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_05850_),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\line_cache[87][1] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_04540_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\line_cache[166][5] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_06071_),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\line_cache[109][2] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_04945_),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\line_cache[89][5] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_04887_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_04586_),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\line_cache[134][7] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_05454_),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\line_cache[190][7] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_06512_),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\line_cache[189][6] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_06492_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\line_cache[173][4] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_06195_),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\line_cache[173][0] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\line_cache[245][4] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_06183_),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\line_cache[166][6] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_06073_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\line_cache[171][0] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_06150_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\line_cache[247][4] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_07548_),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\line_cache[149][1] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_05744_),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\line_cache[261][3] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_07511_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_07806_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\line_cache[261][1] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_07799_),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\line_cache[221][2] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_07070_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\line_cache[94][0] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_04670_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\line_cache[250][6] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_07609_),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\line_cache[150][5] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\line_cache[141][7] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_05776_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\line_cache[143][7] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_05650_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\line_cache[259][4] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_07772_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\line_cache[155][5] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_05866_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\line_cache[169][5] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_06125_),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\line_cache[134][0] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\line_cache[78][7] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_05616_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_05439_),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\line_cache[73][4] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_04288_),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\line_cache[246][2] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_07528_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\line_cache[134][1] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_05441_),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\line_cache[222][2] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_07092_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\line_cache[101][1] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\line_cache[73][0] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_04795_),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\line_cache[74][1] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_04302_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\line_cache[11][6] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_03129_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\line_cache[155][4] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_05864_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\line_cache[165][2] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_06042_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\line_cache[149][3] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_04275_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_05751_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\line_cache[189][1] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_06476_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\line_cache[9][6] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_03094_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\line_cache[270][4] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_07975_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\line_cache[266][4] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_07903_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\line_cache[165][5] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\line_cache[259][5] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_06051_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\line_cache[125][7] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_05283_),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\line_cache[86][6] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_04534_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\line_cache[79][1] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_04394_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\line_cache[86][5] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_04532_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\line_cache[138][1] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_07774_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_05526_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\line_cache[9][2] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_03082_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\line_cache[269][2] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_07949_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\line_cache[74][5] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_04310_),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\line_cache[270][7] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_07981_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\line_cache[239][3] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\line_cache[106][3] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_07399_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\line_cache[189][7] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_06495_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\line_cache[14][6] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_03187_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\line_cache[238][0] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_07376_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\line_cache[239][4] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_07401_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\line_cache[262][2] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_04896_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_07825_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\line_cache[13][3] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_03160_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\line_cache[79][6] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_04404_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\line_cache[149][4] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_05754_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\line_cache[85][6] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_04516_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\line_cache[245][1] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\line_cache[107][1] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_07502_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\line_cache[207][4] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_06822_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\line_cache[153][5] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_05830_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\line_cache[95][4] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_04695_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\line_cache[95][0] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_04686_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\line_cache[242][7] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_04908_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_07464_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\line_cache[91][7] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_04627_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\line_cache[9][0] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_03076_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\line_cache[250][2] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_07601_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\line_cache[270][5] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_07977_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\line_cache[266][3] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\line_cache[69][1] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_07901_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\line_cache[261][2] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_07803_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\line_cache[15][5] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_03202_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\line_cache[126][6] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_05298_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\line_cache[5][2] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_03008_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\line_cache[6][5] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_04390_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_04204_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_03036_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\line_cache[93][6] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_04664_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\line_cache[221][1] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_07066_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\line_cache[111][5] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_04990_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\line_cache[259][2] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_07768_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\line_cache[174][3] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\line_cache[105][3] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_06214_),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\line_cache[205][1] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_06776_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\line_cache[207][0] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_06814_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\line_cache[206][0] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_06797_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\line_cache[85][5] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_04513_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\line_cache[191][5] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_04875_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_06525_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\line_cache[102][1] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_04818_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\line_cache[269][3] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_07952_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\line_cache[269][5] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_07958_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\line_cache[223][4] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_07113_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\line_cache[89][4] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\line_cache[133][2] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_04583_),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\line_cache[102][7] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_04831_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\line_cache[142][0] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_05619_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\line_cache[138][6] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_05541_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\line_cache[71][1] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_04244_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\line_cache[205][7] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_05421_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_06794_),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\line_cache[170][5] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_06144_),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\line_cache[175][5] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_06234_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\line_cache[241][3] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_07435_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\line_cache[191][2] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_06519_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\line_cache[153][4] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\line_cache[77][0] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_05827_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\line_cache[249][5] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_07588_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\line_cache[167][7] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_06091_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\line_cache[257][2] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_07729_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\line_cache[151][2] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_05787_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\line_cache[173][6] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_04351_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_06201_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\line_cache[205][2] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_06779_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\line_cache[171][5] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_06161_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\line_cache[189][3] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_06483_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\line_cache[269][7] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_07964_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\line_cache[110][1] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\line_cache[77][1] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_04965_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\line_cache[95][2] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_04691_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\line_cache[90][4] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_04605_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\line_cache[6][3] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(_03032_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\line_cache[222][0] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(_07088_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\line_cache[265][2] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_04354_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(_07876_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\line_cache[134][6] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_05452_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\line_cache[111][6] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_04992_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\line_cache[126][1] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_05288_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\line_cache[166][1] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_06062_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\line_cache[170][0] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\line_cache[73][3] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_06134_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\line_cache[142][4] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(_05628_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\line_cache[9][7] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(_03097_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\line_cache[238][3] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(_07383_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\line_cache[154][2] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_05844_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\line_cache[74][4] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\line_cache[77][7] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_04285_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(_04308_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\line_cache[6][7] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_03040_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\line_cache[246][7] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_07538_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\line_cache[5][4] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(_03014_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\line_cache[270][3] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(_07973_),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\line_cache[251][7] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\line_cache[241][7] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(_07628_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\line_cache[127][1] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_05304_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\line_cache[75][1] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(_04318_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\line_cache[153][1] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_05818_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\line_cache[250][7] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(_07611_),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\line_cache[238][2] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_07447_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(_07381_),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\line_cache[127][0] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(_05302_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\line_cache[102][6] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_04829_),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\line_cache[191][0] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(_06514_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\line_cache[74][3] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_04306_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\line_cache[151][7] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\line_cache[141][6] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(_05797_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\line_cache[205][5] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(_06788_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\line_cache[239][0] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_07393_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\line_cache[167][2] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_06081_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\line_cache[259][3] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(_07770_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\line_cache[111][4] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_05612_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(_04988_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\line_cache[143][4] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(_05644_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\line_cache[249][4] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(_07585_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\line_cache[237][7] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_07373_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\line_cache[71][4] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_04250_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\line_cache[247][2] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\line_cache[105][4] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(_07544_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\line_cache[77][5] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(_04366_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\line_cache[14][3] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(_03181_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\line_cache[102][5] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(_04827_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\line_cache[75][3] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_04323_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\line_cache[6][6] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_04878_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_03038_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\line_cache[246][6] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_07536_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\line_cache[139][5] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_05563_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\line_cache[243][2] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_07471_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\line_cache[135][5] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_05466_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\line_cache[7][5] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\line_cache[106][5] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(_03053_),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\line_cache[75][0] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_04316_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\line_cache[138][7] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_05544_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\line_cache[102][4] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(_04825_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\line_cache[206][7] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_06812_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\line_cache[150][3] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_04900_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(_05772_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\line_cache[247][1] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(_07542_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\line_cache[221][3] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_07073_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\line_cache[266][0] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_07894_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\line_cache[190][1] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(_06500_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\line_cache[249][3] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\line_cache[125][3] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_07582_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\line_cache[245][2] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(_07505_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\line_cache[155][7] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(_05870_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\line_cache[247][3] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(_07546_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\line_cache[139][4] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_05560_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\line_cache[167][3] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_04372_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_05271_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(_06083_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\line_cache[258][7] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(_07762_),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\line_cache[71][6] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_04254_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\line_cache[222][1] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_07090_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\line_cache[221][6] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_07082_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\line_cache[221][4] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\line_cache[2][0] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_07076_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\line_cache[239][6] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_07405_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\line_cache[6][2] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_03030_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\line_cache[165][3] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_06045_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\line_cache[207][7] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(_06828_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\line_cache[133][6] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_02914_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(_05433_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\line_cache[206][1] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_06799_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\line_cache[71][7] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(_04256_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\line_cache[71][3] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(_04248_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\line_cache[239][1] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(_07395_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\line_cache[238][7] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\line_cache[267][6] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_07391_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\line_cache[222][6] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(_07100_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\line_cache[75][2] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(_04321_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\line_cache[139][2] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_05554_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\line_cache[154][1] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(_05841_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\line_cache[6][0] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_07923_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_03026_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\line_cache[135][2] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(_05460_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\line_cache[149][5] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(_05757_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\line_cache[242][0] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(_07450_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\line_cache[249][2] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_07579_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\line_cache[167][4] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\line_cache[1][4] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(_06085_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\line_cache[3][1] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(_02958_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\line_cache[74][2] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_04304_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\line_cache[270][1] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_07969_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\line_cache[241][5] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(_07441_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\line_cache[102][2] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_02887_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(_04821_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\line_cache[7][0] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(_03042_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\line_cache[7][3] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(_03049_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\line_cache[251][1] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(_07615_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\line_cache[167][5] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(_06087_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\line_cache[205][0] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\line_cache[133][3] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(_06773_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\line_cache[223][5] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_07115_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\pixel_double_counter[3] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_02795_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(_00174_),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\line_cache[85][0] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(_04497_),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\line_cache[251][6] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(_07626_),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_05424_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\line_cache[243][0] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(_07466_),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\line_cache[237][4] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(_07364_),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\line_cache[138][2] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(_05529_),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\line_cache[86][0] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(_04522_),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\line_cache[190][6] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(_06510_),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\line_cache[166][2] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(\line_cache[154][0] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(_05839_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\line_cache[3][5] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(_02974_),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\line_cache[10][6] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(_03113_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\line_cache[71][5] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(_04252_),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\line_cache[15][4] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(_03200_),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\line_cache[105][2] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_06065_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\line_cache[94][5] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(_04680_),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\line_cache[243][1] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(_07468_),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\line_cache[153][2] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(_05821_),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\line_cache[11][4] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(_03125_),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\line_cache[13][0] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(_03150_),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\line_cache[77][6] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\line_cache[269][1] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(_07945_),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\line_cache[158][7] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(_05928_),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\line_cache[251][5] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(_07624_),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\line_cache[247][6] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(_07552_),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\line_cache[15][7] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(_03206_),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_04369_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\line_cache[154][7] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_05854_),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\line_cache[13][1] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(_03153_),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\line_cache[251][0] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(_07613_),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\line_cache[206][3] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(_06804_),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\line_cache[205][3] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(_06782_),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\line_cache[106][0] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\line_cache[159][2] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(_05935_),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(\line_cache[251][2] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(_07618_),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(\line_cache[221][7] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(_07085_),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\line_cache[157][4] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(_05902_),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\line_cache[3][3] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(_02966_),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_04890_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\line_cache[159][4] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(_05939_),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(\line_cache[222][4] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\line_cache[241][2] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_07432_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\line_cache[239][7] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\line_cache[7][1] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(_03044_),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(\line_cache[11][3] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(_03123_),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\line_cache[93][1] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\line_cache[90][0] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\pixel_double_counter[2] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(_02791_),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(_00173_),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(\line_cache[170][2] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\line_cache[15][3] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(_03198_),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\line_cache[250][3] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(_07603_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\line_cache[222][3] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_04648_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_07094_),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\line_cache[3][4] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\line_cache[149][0] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\line_cache[171][2] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\line_cache[158][4] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\line_cache[169][0] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(\line_cache[13][2] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\line_cache[205][6] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_06791_),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\line_cache[149][2] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\line_cache[245][7] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\res_h_counter[9] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(_00160_),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\line_cache[241][6] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\line_cache[3][2] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(\line_cache[207][1] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\line_cache[171][4] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_06159_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\line_cache[170][4] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\line_cache[153][0] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\line_cache[14][0] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_07520_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\line_cache[242][2] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\line_cache[14][1] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(\line_cache[7][4] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\line_cache[222][7] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\line_cache[242][1] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\line_cache[13][7] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(\line_cache[15][0] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\line_cache[14][2] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\line_cache[223][7] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\line_cache[223][6] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\line_cache[261][5] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(\line_cache[133][5] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\line_cache[242][6] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(\line_cache[15][1] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\line_cache[14][5] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\line_cache[13][5] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\line_cache[15][2] ),
    .X(net1984));
 sky130_fd_sc_hd__clkbuf_2 hold1596 (.A(\base_h_counter[0] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(_00131_),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\line_cache[133][1] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\line_cache[251][3] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_04872_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_07812_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(\line_cache[247][7] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\line_cache[14][7] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(\line_cache[251][4] ),
    .X(net1991));
 sky130_fd_sc_hd__buf_1 hold1603 (.A(\line_double_counter[2] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_00177_),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\fb_read_state[0] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_09060_),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(_00009_),
    .X(net1996));
 sky130_fd_sc_hd__clkbuf_2 hold1608 (.A(\res_h_counter[6] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(_00157_),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\line_cache[11][5] ),
    .X(net550));
 sky130_fd_sc_hd__buf_1 hold1610 (.A(\pixel_double_counter[1] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(_02786_),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_00172_),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\line_cache[207][2] ),
    .X(net2002));
 sky130_fd_sc_hd__buf_1 hold1614 (.A(\res_v_counter[1] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(_00162_),
    .X(net2004));
 sky130_fd_sc_hd__buf_1 hold1616 (.A(\line_double_counter[3] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(_00178_),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(net120),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(_00063_),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_03127_),
    .X(net551));
 sky130_fd_sc_hd__buf_1 hold1620 (.A(net110),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(_00053_),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\base_v_counter[2] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(_12878_),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_00143_),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\pixel_double_counter[0] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(_02781_),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(_00171_),
    .X(net2016));
 sky130_fd_sc_hd__buf_1 hold1628 (.A(net118),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_00061_),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\line_cache[133][0] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\line_cache[21][1] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\line_cache[0][1] ),
    .X(net2020));
 sky130_fd_sc_hd__buf_1 hold1632 (.A(net114),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_00057_),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\line_cache[224][4] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\line_cache[181][0] ),
    .X(net2024));
 sky130_fd_sc_hd__buf_1 hold1636 (.A(\base_v_counter[0] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(_12838_),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_00141_),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\res_v_counter[8] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_05415_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_00169_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\line_cache[204][6] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\line_cache[104][1] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\line_cache[244][7] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\line_cache[260][1] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\line_cache[21][7] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\line_cache[183][0] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\line_cache[63][3] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(\line_cache[76][1] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\line_cache[212][2] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\line_cache[223][0] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\line_cache[227][7] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\line_cache[256][2] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\line_cache[244][6] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\line_cache[212][6] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\line_cache[226][2] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\line_cache[128][0] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\line_cache[224][3] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\line_cache[63][2] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(\line_cache[163][1] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\line_cache[240][5] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_07104_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\line_cache[193][5] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\line_cache[0][3] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\line_cache[76][3] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\line_cache[260][3] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\line_cache[192][6] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\line_cache[225][4] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(\line_cache[244][3] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\line_cache[76][0] ),
    .X(net2056));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1668 (.A(\res_v_counter[9] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(_00170_),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\line_cache[103][0] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(\line_cache[63][7] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\line_cache[225][3] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\line_cache[214][7] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\line_cache[228][7] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(\line_cache[212][0] ),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\line_cache[182][4] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\line_cache[214][4] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\line_cache[229][6] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\line_cache[228][3] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\line_cache[182][5] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_04833_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\line_cache[128][7] ),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\line_cache[213][5] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\line_cache[227][4] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\line_cache[227][5] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\line_cache[211][6] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\line_cache[181][5] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\line_cache[192][2] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\line_cache[214][5] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\line_cache[225][7] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\line_cache[182][2] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\line_cache[257][7] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\line_cache[302][1] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\line_cache[302][0] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\line_cache[63][1] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\line_cache[182][6] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\line_cache[244][5] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\line_cache[181][6] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\line_cache[213][6] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\line_cache[76][2] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(\line_cache[211][2] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\line_cache[21][2] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\line_cache[1][7] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_07744_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\line_cache[224][5] ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\line_cache[226][1] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\line_cache[302][5] ),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\line_cache[211][3] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\line_cache[128][2] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\line_cache[302][7] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\line_cache[227][6] ),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\line_cache[225][1] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\line_cache[63][6] ),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\line_cache[181][7] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\line_cache[70][2] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\line_cache[104][6] ),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\line_cache[264][3] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\line_cache[21][5] ),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\line_cache[211][5] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\line_cache[256][7] ),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\line_cache[229][5] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(\line_cache[12][7] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\line_cache[228][0] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(\line_cache[228][4] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\line_cache[182][1] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_04230_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\line_cache[244][2] ),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\line_double_counter[0] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(_02800_),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(_00175_),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\line_cache[21][3] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\line_cache[240][6] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\line_cache[226][6] ),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\line_cache[302][4] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\line_cache[193][6] ),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\line_cache[121][1] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\line_cache[261][0] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\line_cache[244][4] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\line_cache[220][7] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\line_cache[212][3] ),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\line_cache[224][6] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\line_cache[240][4] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(\line_cache[121][4] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\line_cache[212][7] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\line_cache[76][6] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(\line_cache[226][5] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\line_cache[302][6] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_07796_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\line_cache[229][7] ),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\line_cache[42][0] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\line_cache[182][7] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\line_cache[226][0] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\line_cache[302][2] ),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\line_cache[211][7] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(\line_cache[307][2] ),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\line_cache[192][3] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\line_cache[104][3] ),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\line_cache[104][7] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\line_cache[169][7] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\line_cache[181][1] ),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\line_cache[227][1] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\line_cache[213][0] ),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\line_cache[227][0] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\line_cache[163][3] ),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\line_cache[256][6] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\line_cache[213][3] ),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\line_cache[213][4] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\line_cache[193][3] ),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\line_cache[88][2] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_06131_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\line_cache[56][7] ),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\line_cache[313][1] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(\line_cache[260][0] ),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\line_cache[48][0] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\line_cache[244][1] ),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\line_cache[97][7] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(\line_cache[181][4] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\line_cache[236][5] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(\line_cache[12][5] ),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\line_cache[99][1] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\line_cache[258][5] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(\line_cache[278][0] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\line_cache[204][0] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(\line_cache[67][7] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\line_cache[104][5] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\line_cache[200][3] ),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\line_cache[226][3] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(\line_cache[227][3] ),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\line_cache[193][2] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\line_cache[227][2] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\line_cache[41][0] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_07758_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(\line_cache[145][0] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\line_cache[228][2] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\line_cache[51][1] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\line_cache[192][0] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(\line_cache[212][5] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\line_cache[228][1] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(\line_cache[42][2] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\line_cache[81][3] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(\line_cache[183][1] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\line_cache[63][0] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\line_cache[107][7] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(\line_cache[264][5] ),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\line_cache[204][2] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(\line_cache[96][6] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\line_cache[224][1] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(\line_cache[279][4] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\line_cache[121][5] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(\line_cache[38][2] ),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\line_cache[92][7] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(\line_cache[193][0] ),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\line_cache[217][2] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_02908_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_04921_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\line_cache[48][2] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\line_cache[12][1] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(\line_cache[226][7] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\line_cache[4][3] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\line_cache[225][5] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\line_cache[212][1] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\line_cache[104][2] ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\line_cache[179][0] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(\line_cache[208][6] ),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\line_cache[48][1] ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\line_cache[111][1] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(\line_cache[21][6] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\line_cache[260][4] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(\line_cache[156][4] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\line_cache[292][0] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(\line_cache[284][2] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\line_cache[192][1] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(\line_cache[4][7] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\line_cache[152][5] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\line_cache[123][7] ),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\line_cache[37][1] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_04982_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(\line_cache[19][2] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\line_cache[256][3] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(\line_cache[256][5] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\line_cache[244][0] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(\line_cache[59][5] ),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\line_cache[216][6] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(\line_cache[58][4] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(\line_cache[161][2] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(\line_cache[148][4] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(\line_cache[76][7] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\line_cache[133][4] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(\line_cache[161][5] ),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(\line_cache[225][6] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(\line_cache[65][1] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(\line_cache[12][4] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(\line_cache[42][3] ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\line_cache[312][7] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(\line_cache[4][1] ),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\line_cache[216][5] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(\line_cache[296][0] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\line_cache[92][6] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_05427_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(\line_cache[194][7] ),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\line_cache[162][5] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(\line_cache[284][4] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\line_cache[163][6] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(\line_cache[216][2] ),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\line_cache[88][4] ),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(\line_cache[161][6] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(\line_cache[181][2] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(\line_cache[61][1] ),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\line_cache[72][5] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\line_cache[171][3] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(\line_cache[38][0] ),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(\line_cache[305][1] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(\line_cache[16][1] ),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(\line_cache[197][3] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(\line_cache[37][2] ),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(\line_cache[208][3] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(\line_cache[284][5] ),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(\line_cache[51][2] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(\line_cache[292][6] ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(\line_cache[161][1] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_06157_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(\line_cache[296][6] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(\line_cache[4][2] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(\line_cache[252][4] ),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(\line_cache[180][7] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(\line_cache[292][2] ),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(\line_cache[193][4] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(\line_cache[56][1] ),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(\line_cache[163][5] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(\line_cache[182][3] ),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(\line_cache[283][0] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\line_cache[174][2] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(\line_cache[180][0] ),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(\line_cache[0][0] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(\line_cache[308][7] ),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(\line_cache[48][6] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(\line_cache[203][7] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(\line_cache[273][5] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(\line_cache[37][6] ),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(\line_cache[226][4] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(\line_cache[56][4] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(\line_cache[180][1] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_06212_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(\line_cache[28][6] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\line_cache[22][0] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(\line_cache[229][0] ),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(\line_cache[300][5] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(\line_cache[148][3] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(\line_cache[21][4] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(\line_cache[217][1] ),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\line_cache[116][1] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(\line_cache[80][7] ),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(\line_cache[282][3] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\line_cache[125][5] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(\line_cache[288][6] ),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(\line_cache[313][4] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(\line_cache[123][4] ),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(\line_cache[181][3] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(\line_cache[38][4] ),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(\line_cache[256][0] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(\line_cache[163][7] ),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(\line_cache[288][0] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(\line_cache[208][7] ),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(\line_cache[185][2] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\line_cache[78][3] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_05277_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(\line_cache[140][3] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(\line_cache[68][3] ),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(\line_cache[63][5] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\line_cache[185][3] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(\line_cache[37][0] ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(\line_cache[316][2] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(\line_cache[192][4] ),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(\line_cache[233][1] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(\line_cache[284][3] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(\line_cache[160][0] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\line_cache[109][1] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(\line_cache[276][4] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(\line_cache[53][1] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(\line_cache[229][3] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(\line_cache[81][5] ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(\line_cache[49][6] ),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(\line_cache[315][7] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(\line_cache[193][7] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(\line_cache[131][6] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(\line_cache[292][7] ),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(\line_cache[301][0] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_04942_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(\line_cache[224][7] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(\line_cache[280][2] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(\line_cache[317][4] ),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(\line_cache[274][7] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(\line_cache[30][1] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(\line_cache[59][6] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(\line_cache[275][3] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(\line_cache[92][0] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(\line_cache[12][2] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(\line_cache[22][6] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\line_cache[245][0] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(\line_cache[65][0] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\line_cache[308][0] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(\line_cache[304][6] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(\line_cache[12][3] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(\line_cache[26][0] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(\line_cache[99][0] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(\line_cache[194][5] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(\line_cache[56][3] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(\line_cache[230][6] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(\line_cache[208][4] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_07499_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(\line_cache[291][4] ),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(\line_cache[298][3] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(\line_cache[180][3] ),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(\line_cache[260][2] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(\line_cache[290][2] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\line_cache[196][2] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(\line_cache[216][3] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(\line_cache[4][6] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(\line_cache[231][7] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(\line_cache[32][2] ),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\line_cache[11][1] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(\line_cache[42][6] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\line_cache[268][3] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(\line_cache[96][1] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(\line_cache[275][7] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(\line_cache[34][5] ),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(\line_cache[256][1] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(\line_cache[32][4] ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(\line_cache[147][0] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(\line_cache[8][2] ),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(\line_cache[0][6] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_03119_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(\line_cache[275][4] ),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(\line_cache[288][4] ),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(\line_cache[18][3] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(\line_cache[60][3] ),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(\line_cache[188][0] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(\line_cache[211][0] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(\line_cache[236][1] ),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(\line_cache[22][2] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(\line_cache[115][4] ),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(\line_cache[41][1] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\line_cache[109][4] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(\line_cache[33][0] ),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(\line_cache[299][6] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(\line_cache[21][0] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(\line_cache[0][2] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(\line_cache[252][1] ),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(\line_cache[81][1] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(\line_cache[161][0] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(\line_cache[147][4] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(\line_cache[240][7] ),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(\line_cache[84][3] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_04951_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(\line_cache[152][6] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(\line_cache[63][4] ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(\line_cache[41][7] ),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(\line_cache[65][6] ),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(\line_cache[309][5] ),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(\line_cache[8][6] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(\line_cache[240][0] ),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(\line_cache[54][0] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(\line_cache[41][6] ),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(\line_cache[214][0] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\line_cache[243][7] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(\line_cache[119][3] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(\line_cache[278][7] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(\line_cache[193][1] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\line_cache[99][3] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(\line_cache[49][2] ),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(\line_cache[88][6] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(\line_cache[304][0] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(\line_cache[311][1] ),
    .X(net2386));
 sky130_fd_sc_hd__buf_1 hold1998 (.A(net4004),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(\line_cache[49][0] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_04884_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_04382_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_07481_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(\line_cache[62][6] ),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(\line_cache[314][1] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(\line_cache[200][4] ),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(\line_cache[186][1] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(\line_cache[117][0] ),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(\line_cache[281][2] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(\line_cache[114][7] ),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(\line_cache[232][0] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(\line_cache[176][6] ),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(\line_cache[53][7] ),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\line_cache[262][0] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(\line_cache[230][1] ),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(\line_cache[45][3] ),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(\line_cache[120][2] ),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(\line_cache[194][0] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(\line_cache[248][7] ),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(\line_cache[45][4] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(\line_cache[26][7] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(\line_cache[50][2] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(\line_cache[199][3] ),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(\line_cache[209][3] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_07821_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(\line_cache[230][7] ),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(\line_cache[147][2] ),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(\line_cache[231][4] ),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(\line_cache[300][4] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(\line_cache[83][3] ),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(\line_cache[51][5] ),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(\line_cache[26][2] ),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(\line_cache[46][5] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(\line_cache[16][2] ),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(\line_cache[201][7] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\line_cache[107][4] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(\line_cache[197][0] ),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(\line_cache[148][1] ),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(\line_cache[280][7] ),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(\line_cache[299][4] ),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(\line_cache[197][7] ),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(\line_cache[309][4] ),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(\line_cache[97][0] ),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(\line_cache[199][0] ),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(\line_cache[187][4] ),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(\line_cache[81][6] ),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_04915_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(\line_cache[280][0] ),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(\line_cache[273][6] ),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(\line_cache[148][5] ),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(\line_cache[218][1] ),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(\line_cache[20][2] ),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(\line_cache[304][3] ),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(\line_cache[214][6] ),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(\line_cache[218][3] ),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(\line_cache[104][0] ),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(\line_cache[62][1] ),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\line_cache[242][4] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(\line_cache[281][4] ),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(\line_cache[38][1] ),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2052 (.A(\line_cache[113][2] ),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(\line_cache[231][0] ),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(\line_cache[177][2] ),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(\line_cache[275][2] ),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(\line_cache[45][0] ),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(\line_cache[59][0] ),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(\line_cache[240][3] ),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(\line_cache[46][3] ),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_07458_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2060 (.A(\line_cache[295][6] ),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(\line_cache[312][3] ),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2062 (.A(\line_cache[41][2] ),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(\line_cache[302][3] ),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(\line_cache[29][6] ),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(\line_cache[27][0] ),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2066 (.A(\line_cache[97][3] ),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(\line_cache[50][5] ),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(\line_cache[217][3] ),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(\line_cache[177][1] ),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\line_cache[10][1] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(\line_cache[296][3] ),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2071 (.A(\line_cache[46][6] ),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(\line_cache[47][6] ),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(\line_cache[37][4] ),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(\line_cache[148][7] ),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(\line_cache[130][3] ),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2076 (.A(\line_cache[185][0] ),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2077 (.A(\line_cache[177][5] ),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(\line_cache[82][0] ),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(\line_cache[36][1] ),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_03102_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(\line_cache[310][4] ),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2081 (.A(\line_cache[196][7] ),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(\line_cache[288][2] ),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(\line_cache[115][3] ),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(\line_cache[50][1] ),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(\line_cache[17][5] ),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(\line_cache[231][3] ),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2087 (.A(\line_cache[80][2] ),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2088 (.A(\line_cache[28][5] ),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(\line_cache[292][1] ),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\line_cache[271][6] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(\line_cache[297][5] ),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(\line_cache[283][7] ),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(\line_cache[277][3] ),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(\line_cache[230][5] ),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(\line_cache[291][7] ),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(\line_cache[312][4] ),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(\line_cache[202][2] ),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2097 (.A(\line_cache[26][6] ),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(\line_cache[305][4] ),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(\line_cache[162][7] ),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\line_cache[78][2] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_07995_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(\line_cache[72][1] ),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2101 (.A(\line_cache[298][6] ),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(\line_cache[273][2] ),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(\line_cache[52][6] ),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(\line_cache[284][0] ),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2105 (.A(\line_cache[56][5] ),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(\line_cache[68][5] ),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(\line_cache[54][7] ),
    .X(net2496));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2108 (.A(\res_v_counter[4] ),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(_00165_),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\line_cache[109][7] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(\line_cache[37][5] ),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(\line_cache[301][3] ),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2112 (.A(\line_cache[18][7] ),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(\line_cache[276][6] ),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(\line_cache[278][2] ),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(\line_cache[252][0] ),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2116 (.A(\line_cache[160][2] ),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2117 (.A(\line_cache[200][7] ),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(\line_cache[40][2] ),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(\line_cache[234][5] ),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_04960_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(\line_cache[278][4] ),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(\line_cache[184][2] ),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2122 (.A(\line_cache[276][0] ),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2123 (.A(\line_cache[114][4] ),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(\line_cache[25][5] ),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(\line_cache[216][4] ),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(\line_cache[314][7] ),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2127 (.A(\line_cache[291][6] ),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2128 (.A(\line_cache[313][7] ),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(\line_cache[306][0] ),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\line_cache[107][2] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(\line_cache[124][1] ),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(\line_cache[128][1] ),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(\line_cache[140][1] ),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2133 (.A(\line_cache[97][5] ),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(\line_cache[184][0] ),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(\line_cache[25][0] ),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(\line_cache[192][5] ),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(\line_cache[273][7] ),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(\line_cache[299][2] ),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2139 (.A(\line_cache[80][1] ),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_04911_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(\line_cache[214][3] ),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(\line_cache[64][7] ),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(\line_cache[23][0] ),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(\line_cache[192][7] ),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(\line_cache[45][7] ),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2145 (.A(\line_cache[313][3] ),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(\line_cache[72][3] ),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(\line_cache[26][1] ),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(\line_cache[187][2] ),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(\line_cache[51][3] ),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\line_cache[70][1] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(\line_cache[161][4] ),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2151 (.A(\line_cache[216][1] ),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(\line_cache[307][1] ),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2153 (.A(\line_cache[280][4] ),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(\line_cache[26][4] ),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(\line_cache[306][3] ),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(\line_cache[64][3] ),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2157 (.A(\line_cache[46][2] ),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2158 (.A(\line_cache[132][3] ),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(\line_cache[96][7] ),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_04227_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(\line_cache[100][1] ),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(\line_cache[264][0] ),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2162 (.A(\line_cache[295][0] ),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(\line_cache[202][3] ),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(\line_cache[295][7] ),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(\line_cache[299][5] ),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(\line_cache[295][2] ),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(\line_cache[279][2] ),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(\line_cache[117][1] ),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2169 (.A(\line_cache[310][1] ),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\line_cache[190][4] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(\line_cache[220][4] ),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(\line_cache[22][5] ),
    .X(net2560));
 sky130_fd_sc_hd__buf_1 hold2172 (.A(net93),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2173 (.A(_00036_),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(\line_cache[279][1] ),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(\line_cache[182][0] ),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(\line_cache[172][5] ),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(\line_cache[132][5] ),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(\line_cache[293][7] ),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2179 (.A(\line_cache[218][4] ),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_06506_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(\line_cache[307][3] ),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2181 (.A(\line_cache[33][2] ),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(\line_cache[307][7] ),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(\line_cache[309][1] ),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2184 (.A(\line_cache[60][1] ),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(\line_cache[186][5] ),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(\line_cache[128][6] ),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(\line_cache[315][2] ),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(\line_cache[60][5] ),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2189 (.A(\line_cache[303][2] ),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\line_cache[2][7] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(\line_cache[315][4] ),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2191 (.A(\line_cache[285][5] ),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(\line_cache[108][7] ),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(\line_cache[188][6] ),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(\line_cache[42][5] ),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(\line_cache[232][1] ),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(\line_cache[278][5] ),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2197 (.A(\line_cache[188][3] ),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(\line_cache[144][4] ),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2199 (.A(\line_cache[55][0] ),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_04380_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_02950_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(\line_cache[129][5] ),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(\line_cache[297][1] ),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2202 (.A(\line_cache[276][1] ),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(\line_cache[220][5] ),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(\line_cache[146][5] ),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(\line_cache[59][3] ),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(\line_cache[131][4] ),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(\line_cache[42][4] ),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(\line_cache[303][6] ),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(\line_cache[314][3] ),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\line_cache[259][0] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(\line_cache[217][0] ),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(\line_cache[68][7] ),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(\line_cache[35][1] ),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(\line_cache[176][5] ),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(\line_cache[160][4] ),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2215 (.A(\line_cache[27][3] ),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(\line_cache[277][2] ),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(\line_cache[19][1] ),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(\line_cache[45][1] ),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(\line_cache[285][4] ),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_07764_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(\line_cache[81][2] ),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(\line_cache[65][2] ),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(\line_cache[19][3] ),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(\line_cache[23][2] ),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(\line_cache[272][6] ),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(\line_cache[55][3] ),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(\line_cache[195][2] ),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2227 (.A(\line_cache[303][3] ),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(\line_cache[152][1] ),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(\line_cache[308][2] ),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\line_cache[86][2] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(\line_cache[160][7] ),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(\line_cache[23][3] ),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2232 (.A(\line_cache[288][1] ),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(\line_cache[28][0] ),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(\line_cache[311][3] ),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(\line_cache[309][0] ),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(\line_cache[303][5] ),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2237 (.A(\line_cache[304][7] ),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(\line_cache[216][0] ),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(\line_cache[47][1] ),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_04526_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(\line_cache[188][7] ),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(\line_cache[274][6] ),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2242 (.A(\line_cache[232][3] ),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2243 (.A(\line_cache[290][7] ),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2244 (.A(\line_cache[45][2] ),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2245 (.A(\line_cache[104][4] ),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(\line_cache[144][3] ),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(\line_cache[236][6] ),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(\line_cache[81][4] ),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2249 (.A(\line_cache[218][7] ),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\line_cache[86][1] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2250 (.A(\line_cache[152][4] ),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(\line_cache[289][5] ),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2252 (.A(\line_cache[252][2] ),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(\line_cache[200][5] ),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2254 (.A(\line_cache[26][5] ),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(\line_cache[307][4] ),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(\line_cache[229][1] ),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(\line_cache[297][6] ),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(\line_cache[231][2] ),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2259 (.A(\line_cache[177][3] ),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_04524_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(\line_cache[18][4] ),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(\line_cache[96][3] ),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2262 (.A(\line_cache[51][6] ),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2263 (.A(\line_cache[233][2] ),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(\line_cache[185][6] ),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2265 (.A(\line_cache[33][1] ),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(\line_cache[283][5] ),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2267 (.A(\line_cache[66][1] ),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(\line_cache[291][0] ),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(\line_cache[129][7] ),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\line_cache[267][2] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(\line_cache[180][2] ),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2271 (.A(\line_cache[314][4] ),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(\line_cache[131][2] ),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(\line_cache[50][6] ),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2274 (.A(\line_cache[100][0] ),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(\line_cache[62][7] ),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2276 (.A(\line_cache[289][0] ),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(\line_cache[296][2] ),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2278 (.A(\line_cache[314][5] ),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2279 (.A(\line_cache[212][4] ),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_07915_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(\line_cache[194][4] ),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2281 (.A(\line_cache[316][7] ),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(\line_cache[38][5] ),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2283 (.A(\line_cache[34][0] ),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2284 (.A(\line_cache[178][3] ),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2285 (.A(\line_cache[276][5] ),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(\line_cache[156][0] ),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(\line_cache[8][3] ),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(\line_cache[16][7] ),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2289 (.A(\line_cache[301][4] ),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\line_cache[246][0] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(\line_cache[41][4] ),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(\line_cache[268][1] ),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(\line_cache[299][0] ),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(\line_cache[196][4] ),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(\line_cache[194][2] ),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(\line_cache[124][6] ),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(\line_cache[108][2] ),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(\line_cache[8][0] ),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(\line_cache[29][4] ),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2299 (.A(\line_cache[131][5] ),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\line_cache[78][4] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_07523_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2300 (.A(\line_cache[274][0] ),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2301 (.A(\line_cache[64][1] ),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(\line_cache[316][1] ),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(\line_cache[273][4] ),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(\line_cache[17][6] ),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(\line_cache[307][5] ),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2306 (.A(\line_cache[164][4] ),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2307 (.A(\line_cache[68][6] ),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(\line_cache[99][2] ),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(\line_cache[303][0] ),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\line_cache[89][2] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2310 (.A(\line_cache[201][4] ),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(\line_cache[51][4] ),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2312 (.A(\line_cache[161][3] ),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2313 (.A(\line_cache[88][1] ),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(\line_cache[61][3] ),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2315 (.A(\line_cache[146][0] ),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(\line_cache[186][3] ),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(\line_cache[297][3] ),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2318 (.A(\line_cache[53][0] ),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2319 (.A(\line_cache[30][3] ),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_04577_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(\line_cache[311][6] ),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2321 (.A(\line_cache[213][7] ),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2322 (.A(\line_cache[281][7] ),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(\line_cache[196][6] ),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2324 (.A(\line_cache[12][0] ),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(\line_cache[183][4] ),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2326 (.A(\line_cache[152][7] ),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(\line_cache[209][2] ),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(\line_cache[123][2] ),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(\line_cache[308][5] ),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\line_cache[175][6] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(\line_cache[114][2] ),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2331 (.A(\line_cache[50][7] ),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(\line_cache[185][7] ),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2333 (.A(\line_cache[274][5] ),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(\line_cache[35][4] ),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(\line_cache[240][2] ),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2336 (.A(\line_cache[66][0] ),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(\line_cache[27][1] ),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2338 (.A(\line_cache[72][7] ),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(\line_cache[301][6] ),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_06236_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2340 (.A(\line_cache[198][3] ),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(\line_cache[311][2] ),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2342 (.A(\line_cache[4][0] ),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2343 (.A(\line_cache[187][3] ),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2344 (.A(\line_cache[16][6] ),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2345 (.A(\line_cache[62][4] ),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2346 (.A(\line_cache[25][7] ),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2347 (.A(\line_cache[27][4] ),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(\line_cache[65][4] ),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(\line_cache[100][5] ),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\line_cache[11][2] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(\line_cache[294][5] ),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2351 (.A(\line_cache[313][2] ),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2352 (.A(\line_cache[199][2] ),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(\line_cache[294][6] ),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2354 (.A(\line_cache[81][7] ),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2355 (.A(\line_cache[56][2] ),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(\line_cache[66][5] ),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(\line_cache[233][3] ),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(\line_cache[118][4] ),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(\line_cache[196][3] ),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_03121_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2360 (.A(\line_cache[98][0] ),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(net100),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2362 (.A(_00043_),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2363 (.A(\line_cache[61][2] ),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2364 (.A(\line_cache[76][5] ),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(\line_cache[18][0] ),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(\line_cache[58][5] ),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(\line_cache[225][2] ),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(\line_cache[297][4] ),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2369 (.A(\line_cache[306][1] ),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\line_cache[159][6] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2370 (.A(\line_cache[119][1] ),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2371 (.A(\line_cache[234][4] ),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2372 (.A(\line_cache[68][0] ),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(\line_cache[290][1] ),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2374 (.A(\line_cache[16][3] ),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2375 (.A(\line_cache[272][1] ),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2376 (.A(\line_cache[26][3] ),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(\line_cache[313][6] ),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2378 (.A(\line_cache[200][1] ),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2379 (.A(\line_cache[38][3] ),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_05943_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(\line_cache[56][6] ),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2381 (.A(\line_cache[168][3] ),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2382 (.A(\line_cache[35][7] ),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2383 (.A(\line_cache[4][5] ),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(\line_cache[236][0] ),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2385 (.A(\line_cache[300][3] ),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(\line_cache[19][4] ),
    .X(net2775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2387 (.A(\line_cache[18][5] ),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2388 (.A(\line_cache[234][2] ),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(\line_cache[172][4] ),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\line_cache[245][6] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2390 (.A(\line_cache[97][6] ),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2391 (.A(\line_cache[124][2] ),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(\line_cache[23][1] ),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2393 (.A(\line_cache[196][0] ),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2394 (.A(\line_cache[49][5] ),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(\line_cache[180][5] ),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2396 (.A(\line_cache[168][4] ),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(\line_cache[296][5] ),
    .X(net2786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(\line_cache[277][4] ),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(\line_cache[147][7] ),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_04384_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_07517_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2400 (.A(\line_cache[140][0] ),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2401 (.A(\line_cache[119][5] ),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2402 (.A(\line_cache[308][3] ),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2403 (.A(\line_cache[147][3] ),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(\line_cache[35][2] ),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(\line_cache[108][0] ),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2406 (.A(\line_cache[145][1] ),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2407 (.A(\line_cache[29][0] ),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(\line_double_counter[1] ),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(_00176_),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\line_cache[85][2] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(\line_cache[36][2] ),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2411 (.A(\line_cache[33][6] ),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2412 (.A(\line_cache[177][4] ),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(\line_cache[317][0] ),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(\line_cache[140][4] ),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(\line_cache[156][6] ),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2416 (.A(\line_cache[289][2] ),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2417 (.A(\line_cache[38][7] ),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2418 (.A(\line_cache[124][5] ),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(\line_cache[92][1] ),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_04504_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2420 (.A(\line_cache[82][7] ),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(\line_cache[194][3] ),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(\line_cache[29][2] ),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(\line_cache[35][3] ),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2424 (.A(\line_cache[22][7] ),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2425 (.A(\line_cache[114][3] ),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2426 (.A(\line_cache[98][5] ),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(\line_cache[50][4] ),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2428 (.A(\line_cache[275][0] ),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(\line_cache[29][7] ),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\line_cache[267][1] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2430 (.A(\line_cache[232][6] ),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2431 (.A(\line_cache[209][1] ),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2432 (.A(\line_cache[306][5] ),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(\line_cache[186][4] ),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(\line_cache[275][5] ),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(\line_cache[37][7] ),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(\line_cache[37][3] ),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(\line_cache[148][6] ),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(\line_cache[310][7] ),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2439 (.A(\line_cache[23][5] ),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_07913_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(\line_cache[144][7] ),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2441 (.A(\line_cache[30][6] ),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2442 (.A(\line_cache[220][0] ),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(\line_cache[308][4] ),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2444 (.A(\line_cache[129][0] ),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(\line_cache[231][6] ),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(\line_cache[168][1] ),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(\line_cache[60][2] ),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(\line_cache[145][5] ),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(\line_cache[121][3] ),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\line_cache[190][0] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2450 (.A(\line_cache[185][1] ),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2451 (.A(\line_cache[188][2] ),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(\line_cache[234][3] ),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(\line_cache[19][7] ),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2454 (.A(\line_cache[49][3] ),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2455 (.A(\line_cache[96][4] ),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(\line_cache[144][0] ),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(\line_cache[120][1] ),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2458 (.A(\line_cache[156][2] ),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(\line_cache[33][7] ),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_06498_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(\line_cache[315][0] ),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(\line_cache[275][6] ),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2462 (.A(\line_cache[280][1] ),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2463 (.A(\line_cache[168][7] ),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2464 (.A(\line_cache[272][5] ),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(\line_cache[65][3] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(\line_cache[201][1] ),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(\line_cache[117][4] ),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2468 (.A(\line_cache[293][3] ),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2469 (.A(\line_cache[52][7] ),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\line_cache[74][6] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(\line_cache[80][0] ),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2471 (.A(\line_cache[36][0] ),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2472 (.A(\line_cache[209][6] ),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2473 (.A(\line_cache[25][2] ),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(\line_cache[292][5] ),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2475 (.A(\line_cache[112][2] ),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2476 (.A(\line_cache[315][5] ),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(\line_cache[317][3] ),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(\line_cache[209][7] ),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2479 (.A(\line_cache[131][7] ),
    .X(net2868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_04312_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2480 (.A(\line_cache[115][5] ),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(\line_cache[65][7] ),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(\line_cache[317][6] ),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(\line_cache[317][5] ),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2484 (.A(\line_cache[56][0] ),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2485 (.A(\line_cache[231][5] ),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(\line_cache[197][2] ),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2487 (.A(\line_cache[299][3] ),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(\line_cache[283][3] ),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(\line_cache[310][3] ),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\line_cache[73][6] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2490 (.A(\line_cache[316][0] ),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(\line_cache[30][4] ),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2492 (.A(\line_cache[289][3] ),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(\line_cache[60][0] ),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2494 (.A(\line_cache[32][1] ),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(\line_cache[298][7] ),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(\line_cache[272][0] ),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2497 (.A(\line_cache[122][2] ),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2498 (.A(\line_cache[0][7] ),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2499 (.A(\line_cache[228][6] ),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\line_cache[2][4] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_04294_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2500 (.A(\line_cache[291][5] ),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2501 (.A(\line_cache[297][0] ),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2502 (.A(\line_cache[29][5] ),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(\line_cache[307][6] ),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2504 (.A(\line_cache[113][7] ),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2505 (.A(\line_cache[53][4] ),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2506 (.A(\line_cache[147][6] ),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(\line_cache[129][1] ),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2508 (.A(\line_cache[55][6] ),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2509 (.A(\line_cache[8][7] ),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\line_cache[11][0] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2510 (.A(\line_cache[124][3] ),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(\line_cache[88][0] ),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(\line_cache[30][0] ),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(\line_cache[225][0] ),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2514 (.A(\line_cache[136][2] ),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2515 (.A(\line_cache[316][5] ),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2516 (.A(\line_cache[66][2] ),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2517 (.A(\line_cache[168][5] ),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(\line_cache[195][5] ),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2519 (.A(\line_cache[99][5] ),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_03117_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(\line_cache[27][2] ),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2521 (.A(\line_cache[39][2] ),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(\line_cache[30][5] ),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2523 (.A(\line_cache[0][5] ),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(\line_cache[179][3] ),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2525 (.A(\line_cache[279][0] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2526 (.A(\line_cache[301][5] ),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(\line_cache[260][5] ),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2528 (.A(\line_cache[248][4] ),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2529 (.A(\line_cache[64][0] ),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\line_cache[93][2] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2530 (.A(\line_cache[33][3] ),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(\line_cache[22][1] ),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(\line_cache[19][0] ),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(\line_cache[194][6] ),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2534 (.A(\line_cache[42][1] ),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2535 (.A(\line_cache[24][0] ),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(\line_cache[289][6] ),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2537 (.A(\line_cache[23][6] ),
    .X(net2926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2538 (.A(\line_cache[310][0] ),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(\line_cache[28][3] ),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_04652_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2540 (.A(\line_cache[36][4] ),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2541 (.A(\line_cache[146][6] ),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2542 (.A(\line_cache[59][7] ),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(\line_cache[200][6] ),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2544 (.A(\line_cache[54][1] ),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(\line_cache[123][1] ),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2546 (.A(\line_cache[295][1] ),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(\line_cache[252][6] ),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2548 (.A(\line_cache[145][3] ),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(\line_cache[309][6] ),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\line_cache[167][6] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2550 (.A(\line_cache[8][1] ),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2551 (.A(\line_cache[120][3] ),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2552 (.A(\line_cache[232][5] ),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2553 (.A(\line_cache[114][0] ),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(\line_cache[8][4] ),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2555 (.A(\line_cache[268][2] ),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(\line_cache[284][1] ),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2557 (.A(\line_cache[49][4] ),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(\line_cache[217][4] ),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2559 (.A(\line_cache[233][0] ),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_06089_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2560 (.A(\line_cache[252][7] ),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2561 (.A(\line_cache[291][2] ),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2562 (.A(\line_cache[210][5] ),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(\line_cache[289][4] ),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2564 (.A(\line_cache[54][6] ),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2565 (.A(\line_cache[307][0] ),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2566 (.A(\line_cache[294][3] ),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2567 (.A(\line_cache[27][6] ),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2568 (.A(\line_cache[273][1] ),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2569 (.A(\line_cache[66][7] ),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\line_cache[10][2] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2570 (.A(\line_cache[253][0] ),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2571 (.A(\line_cache[84][6] ),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2572 (.A(\line_cache[129][6] ),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2573 (.A(\line_cache[123][3] ),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(\line_cache[80][4] ),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(\line_cache[278][1] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2576 (.A(\line_cache[24][2] ),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2577 (.A(\line_cache[52][4] ),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2578 (.A(\line_cache[285][0] ),
    .X(net2967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(\line_cache[288][5] ),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_03105_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(\line_cache[180][4] ),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(\line_cache[279][3] ),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2582 (.A(\line_cache[116][4] ),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(\line_cache[156][1] ),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(\line_cache[28][1] ),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2585 (.A(\line_cache[311][7] ),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2586 (.A(\line_cache[115][2] ),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(\line_cache[279][6] ),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2588 (.A(\line_cache[116][2] ),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(\line_cache[282][1] ),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\line_cache[159][3] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2590 (.A(\line_cache[289][1] ),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2591 (.A(\line_cache[136][7] ),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(\line_cache[140][6] ),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2593 (.A(\line_cache[48][5] ),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(\line_cache[297][2] ),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(\line_cache[293][4] ),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(\line_cache[81][0] ),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2597 (.A(\line_cache[123][0] ),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2598 (.A(\line_cache[176][1] ),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(\line_cache[84][4] ),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_02935_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_05937_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2600 (.A(\line_cache[64][4] ),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2601 (.A(\line_cache[130][6] ),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2602 (.A(\line_cache[8][5] ),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(\line_cache[178][0] ),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(\line_cache[233][7] ),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2605 (.A(\line_cache[310][2] ),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(\line_cache[268][4] ),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2607 (.A(\line_cache[108][5] ),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(\line_cache[59][4] ),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2609 (.A(\line_cache[289][7] ),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\line_cache[159][5] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2610 (.A(\line_cache[160][1] ),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2611 (.A(\line_cache[195][0] ),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(\line_cache[55][5] ),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(\line_cache[290][5] ),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2614 (.A(\line_cache[60][7] ),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(\line_cache[20][4] ),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(\line_cache[314][0] ),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2617 (.A(\line_cache[220][1] ),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(\line_cache[60][4] ),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(\line_cache[67][0] ),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_05941_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(\line_cache[178][7] ),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2621 (.A(\line_cache[29][1] ),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(\line_cache[292][4] ),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2623 (.A(\line_cache[211][4] ),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2624 (.A(\line_cache[113][5] ),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(\line_cache[41][3] ),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2626 (.A(\line_cache[22][4] ),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2627 (.A(net112),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2628 (.A(_00055_),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(\line_cache[32][3] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\line_cache[95][6] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(\line_cache[123][5] ),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(\line_cache[57][5] ),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2632 (.A(\line_cache[215][7] ),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(\line_cache[312][2] ),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2634 (.A(\line_cache[199][7] ),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(\line_cache[298][2] ),
    .X(net3024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2636 (.A(\line_cache[315][6] ),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2637 (.A(\line_cache[92][4] ),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2638 (.A(\line_cache[17][7] ),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(\line_cache[314][6] ),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_04699_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(\line_cache[301][1] ),
    .X(net3029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2641 (.A(\line_cache[124][4] ),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2642 (.A(\line_cache[184][4] ),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(\line_cache[121][7] ),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(\line_cache[115][1] ),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(\line_cache[136][3] ),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2646 (.A(\line_cache[195][7] ),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2647 (.A(\line_cache[88][7] ),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2648 (.A(\line_cache[313][0] ),
    .X(net3037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(\line_cache[58][7] ),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\line_cache[93][4] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2650 (.A(\line_cache[55][2] ),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(\line_cache[62][3] ),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(\line_cache[33][5] ),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2653 (.A(\line_cache[276][7] ),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(\line_cache[177][7] ),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(\line_cache[100][4] ),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(\line_cache[124][0] ),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(\line_cache[60][6] ),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(\line_cache[311][4] ),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2659 (.A(\line_cache[228][5] ),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_04658_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2660 (.A(\line_cache[20][6] ),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(\line_cache[300][1] ),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2662 (.A(\line_cache[50][0] ),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2663 (.A(\line_cache[122][5] ),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(\line_cache[121][6] ),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2665 (.A(\line_cache[252][3] ),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(\line_cache[232][4] ),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(\line_cache[199][6] ),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(\line_cache[168][2] ),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(\line_cache[117][6] ),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\line_cache[159][0] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(\line_cache[311][5] ),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(\line_cache[136][6] ),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(\line_cache[146][2] ),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(\line_cache[203][2] ),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(\line_cache[285][3] ),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(\line_cache[274][2] ),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(\line_cache[83][1] ),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(\line_cache[298][0] ),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(\line_cache[128][3] ),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(\line_cache[32][7] ),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_05930_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(\line_cache[132][1] ),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(\line_cache[128][4] ),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2682 (.A(\line_cache[303][7] ),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(\line_cache[316][6] ),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(\line_cache[4][4] ),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2685 (.A(\line_cache[306][2] ),
    .X(net3074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(\line_cache[108][4] ),
    .X(net3075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(\line_cache[162][3] ),
    .X(net3076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(\line_cache[248][3] ),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2689 (.A(\line_cache[201][0] ),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\line_cache[190][5] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2690 (.A(\line_cache[282][6] ),
    .X(net3079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(\line_cache[288][3] ),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2692 (.A(\line_cache[177][6] ),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2693 (.A(\line_cache[35][5] ),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2694 (.A(\line_cache[281][0] ),
    .X(net3083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(\line_cache[118][0] ),
    .X(net3084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(\line_cache[278][3] ),
    .X(net3085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2697 (.A(\line_cache[49][1] ),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2698 (.A(\line_cache[294][7] ),
    .X(net3087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(\line_cache[34][2] ),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\line_cache[257][4] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_06508_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(\line_cache[18][6] ),
    .X(net3089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(\line_cache[67][1] ),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(\line_cache[264][7] ),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(\line_cache[278][6] ),
    .X(net3092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(\line_cache[145][4] ),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(\line_cache[305][5] ),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(\line_cache[208][2] ),
    .X(net3095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(\line_cache[279][7] ),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(\line_cache[235][0] ),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2709 (.A(\line_cache[112][7] ),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\line_cache[175][7] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2710 (.A(\line_cache[48][3] ),
    .X(net3099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2711 (.A(\line_cache[49][7] ),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(\line_cache[146][7] ),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2713 (.A(\line_cache[195][6] ),
    .X(net3102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(\line_cache[236][3] ),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(\line_cache[294][1] ),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2716 (.A(\line_cache[290][4] ),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2717 (.A(\line_cache[201][5] ),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2718 (.A(\line_cache[283][4] ),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(\line_cache[32][6] ),
    .X(net3108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_06238_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(\line_cache[184][3] ),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(\line_cache[112][0] ),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2722 (.A(\line_cache[305][3] ),
    .X(net3111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(\line_cache[82][3] ),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(\line_cache[84][0] ),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2725 (.A(\line_cache[219][5] ),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2726 (.A(\line_cache[62][2] ),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(\line_cache[296][1] ),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(\line_cache[130][1] ),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(\line_cache[66][3] ),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\line_cache[87][5] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2730 (.A(\line_cache[98][3] ),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(\line_cache[121][0] ),
    .X(net3120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2732 (.A(\line_cache[129][2] ),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2733 (.A(\line_cache[65][5] ),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2734 (.A(\line_cache[277][5] ),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(\line_cache[113][6] ),
    .X(net3124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(\line_cache[82][2] ),
    .X(net3125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(\line_cache[36][5] ),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2738 (.A(\line_cache[318][3] ),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(\line_cache[52][0] ),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_04549_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2740 (.A(\line_cache[42][7] ),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2741 (.A(\line_cache[100][3] ),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(\line_cache[284][7] ),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(\line_cache[215][0] ),
    .X(net3132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(\line_cache[310][5] ),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(\line_cache[236][7] ),
    .X(net3134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(\line_cache[46][7] ),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(\line_cache[273][3] ),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(\line_cache[180][6] ),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2749 (.A(\line_cache[240][1] ),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\line_cache[261][4] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2750 (.A(\line_cache[234][6] ),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(\line_cache[196][1] ),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2752 (.A(\line_cache[51][0] ),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(\line_cache[296][4] ),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(\line_cache[210][7] ),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2755 (.A(\line_cache[57][3] ),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(\line_cache[160][3] ),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2757 (.A(\line_cache[260][6] ),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2758 (.A(\line_cache[186][2] ),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(\line_cache[118][5] ),
    .X(net3148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_07809_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2760 (.A(\line_cache[54][5] ),
    .X(net3149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2761 (.A(\line_cache[24][7] ),
    .X(net3150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(\line_cache[146][1] ),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(\line_cache[256][4] ),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(\line_cache[97][2] ),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(\line_cache[298][5] ),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(\line_cache[61][0] ),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(\line_cache[46][4] ),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2768 (.A(\line_cache[54][3] ),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2769 (.A(\line_cache[187][5] ),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\line_cache[110][5] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2770 (.A(\line_cache[254][0] ),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(\line_cache[299][7] ),
    .X(net3160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(\line_cache[291][1] ),
    .X(net3161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(\line_cache[122][0] ),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2774 (.A(\line_cache[210][3] ),
    .X(net3163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(\line_cache[202][7] ),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(\line_cache[114][6] ),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(\line_cache[140][7] ),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2778 (.A(\line_cache[301][2] ),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2779 (.A(\line_cache[317][2] ),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_04974_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2780 (.A(\line_cache[293][6] ),
    .X(net3169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(\line_cache[28][2] ),
    .X(net3170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2782 (.A(\line_cache[300][7] ),
    .X(net3171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(\line_cache[248][0] ),
    .X(net3172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2784 (.A(\line_cache[118][1] ),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(\line_cache[272][2] ),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(\line_cache[113][1] ),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2787 (.A(\line_cache[300][0] ),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2788 (.A(\line_cache[236][2] ),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2789 (.A(\line_cache[179][7] ),
    .X(net3178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\line_cache[137][7] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2790 (.A(\line_cache[208][5] ),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(\line_cache[53][6] ),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2792 (.A(\line_cache[201][3] ),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(\line_cache[282][5] ),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(\line_cache[19][6] ),
    .X(net3183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(\line_cache[82][5] ),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(\line_cache[280][3] ),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2797 (.A(\line_cache[100][7] ),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(\line_cache[36][3] ),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2799 (.A(\line_cache[130][4] ),
    .X(net3188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_07735_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_05519_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2800 (.A(\line_cache[217][5] ),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(\line_cache[282][7] ),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(\line_cache[279][5] ),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2803 (.A(\line_cache[34][4] ),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(\line_cache[80][6] ),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(\line_cache[30][2] ),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(\line_cache[309][7] ),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(\line_cache[112][4] ),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2808 (.A(\line_cache[276][2] ),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2809 (.A(\line_cache[12][6] ),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\line_cache[159][1] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2810 (.A(\line_cache[201][2] ),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(\line_cache[54][2] ),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2812 (.A(\line_cache[315][3] ),
    .X(net3201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2813 (.A(\line_cache[34][3] ),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2814 (.A(\line_cache[35][6] ),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(\line_cache[58][0] ),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(\line_cache[280][6] ),
    .X(net3205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(\line_cache[119][6] ),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(\line_cache[55][4] ),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2819 (.A(\line_cache[24][6] ),
    .X(net3208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_05932_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2820 (.A(\line_cache[122][1] ),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2821 (.A(\line_cache[108][6] ),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(\line_cache[303][4] ),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(\line_cache[18][1] ),
    .X(net3212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(\line_cache[130][0] ),
    .X(net3213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(\line_cache[53][3] ),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(\line_cache[198][5] ),
    .X(net3215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(\line_cache[100][6] ),
    .X(net3216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(\line_cache[119][0] ),
    .X(net3217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(\line_cache[198][7] ),
    .X(net3218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\line_cache[91][5] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(\line_cache[84][2] ),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(\line_cache[229][4] ),
    .X(net3220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2832 (.A(\line_cache[66][6] ),
    .X(net3221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(\line_cache[304][4] ),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(\line_cache[176][7] ),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2835 (.A(\line_cache[123][6] ),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(\line_cache[46][0] ),
    .X(net3225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(\line_cache[161][7] ),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2838 (.A(\line_cache[120][5] ),
    .X(net3227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(\line_cache[116][3] ),
    .X(net3228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_04623_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2840 (.A(\line_cache[99][6] ),
    .X(net3229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(\line_cache[52][5] ),
    .X(net3230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(\line_cache[48][4] ),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(\line_cache[308][6] ),
    .X(net3232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(\line_cache[119][4] ),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2845 (.A(\line_cache[176][4] ),
    .X(net3234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2846 (.A(\line_cache[219][4] ),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2847 (.A(\line_cache[197][1] ),
    .X(net3236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(\line_cache[312][5] ),
    .X(net3237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(\line_cache[195][4] ),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\line_cache[107][0] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(\line_cache[220][6] ),
    .X(net3239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(\line_cache[306][4] ),
    .X(net3240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(\line_cache[41][5] ),
    .X(net3241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(\line_cache[132][4] ),
    .X(net3242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2854 (.A(\line_cache[117][5] ),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(\line_cache[185][4] ),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(\line_cache[117][3] ),
    .X(net3245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2857 (.A(\line_cache[64][6] ),
    .X(net3246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(\line_cache[297][7] ),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2859 (.A(\line_cache[98][7] ),
    .X(net3248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_04906_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(\line_cache[288][7] ),
    .X(net3249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2861 (.A(\line_cache[254][2] ),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2862 (.A(\line_cache[310][6] ),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2863 (.A(\line_cache[195][3] ),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2864 (.A(\line_cache[51][7] ),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2865 (.A(\line_cache[82][1] ),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2866 (.A(\line_cache[164][3] ),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2867 (.A(\line_cache[201][6] ),
    .X(net3256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2868 (.A(\line_cache[293][1] ),
    .X(net3257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2869 (.A(\line_cache[53][5] ),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\line_cache[271][3] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2870 (.A(\line_cache[316][4] ),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2871 (.A(\line_cache[172][1] ),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2872 (.A(\line_cache[283][1] ),
    .X(net3261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2873 (.A(\line_cache[254][7] ),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2874 (.A(\line_cache[185][5] ),
    .X(net3263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2875 (.A(\line_cache[97][1] ),
    .X(net3264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2876 (.A(\line_cache[145][7] ),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2877 (.A(\line_cache[24][5] ),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2878 (.A(\line_cache[88][5] ),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2879 (.A(\line_cache[20][3] ),
    .X(net3268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_07989_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2880 (.A(\line_cache[164][2] ),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2881 (.A(\line_cache[132][0] ),
    .X(net3270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2882 (.A(\line_cache[20][7] ),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2883 (.A(\line_cache[224][0] ),
    .X(net3272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2884 (.A(\line_cache[17][2] ),
    .X(net3273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2885 (.A(\line_cache[28][7] ),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2886 (.A(\line_cache[29][3] ),
    .X(net3275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2887 (.A(\line_cache[211][1] ),
    .X(net3276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2888 (.A(\line_cache[32][5] ),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2889 (.A(\line_cache[117][7] ),
    .X(net3278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\line_cache[69][3] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2890 (.A(\line_cache[273][0] ),
    .X(net3279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2891 (.A(\line_cache[36][7] ),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2892 (.A(\line_cache[306][7] ),
    .X(net3281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2893 (.A(\line_cache[210][6] ),
    .X(net3282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2894 (.A(\line_cache[52][2] ),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2895 (.A(\line_cache[34][7] ),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2896 (.A(\line_cache[34][6] ),
    .X(net3285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2897 (.A(\line_cache[306][6] ),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2898 (.A(\line_cache[198][1] ),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2899 (.A(\line_cache[176][3] ),
    .X(net3288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\line_cache[105][1] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_04210_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2900 (.A(\line_cache[131][0] ),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2901 (.A(\line_cache[96][0] ),
    .X(net3290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2902 (.A(\line_cache[294][0] ),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2903 (.A(\line_cache[272][4] ),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2904 (.A(\line_cache[136][0] ),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2905 (.A(\line_cache[67][6] ),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2906 (.A(\line_cache[285][2] ),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2907 (.A(\line_cache[99][7] ),
    .X(net3296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2908 (.A(\line_cache[140][2] ),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2909 (.A(\line_cache[53][2] ),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\line_cache[141][3] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2910 (.A(\line_cache[177][0] ),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2911 (.A(\line_cache[112][1] ),
    .X(net3300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2912 (.A(\line_cache[96][5] ),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2913 (.A(\line_cache[164][5] ),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2914 (.A(\line_cache[313][5] ),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2915 (.A(\line_cache[58][6] ),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2916 (.A(\line_cache[293][0] ),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2917 (.A(\line_cache[152][3] ),
    .X(net3306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2918 (.A(\line_cache[45][5] ),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2919 (.A(\line_cache[184][7] ),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_05600_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2920 (.A(\line_cache[130][7] ),
    .X(net3309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2921 (.A(\line_cache[282][2] ),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2922 (.A(\line_cache[233][4] ),
    .X(net3311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2923 (.A(\line_cache[253][7] ),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2924 (.A(\line_cache[284][6] ),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2925 (.A(\line_cache[168][6] ),
    .X(net3314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2926 (.A(\line_cache[57][4] ),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2927 (.A(\line_cache[220][3] ),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2928 (.A(\line_cache[19][5] ),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2929 (.A(\line_cache[118][3] ),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\line_cache[101][2] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2930 (.A(\line_cache[303][1] ),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2931 (.A(\line_cache[132][7] ),
    .X(net3320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2932 (.A(\line_cache[187][1] ),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2933 (.A(\line_cache[36][6] ),
    .X(net3322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2934 (.A(\line_cache[216][7] ),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2935 (.A(\line_cache[164][7] ),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2936 (.A(\line_cache[144][1] ),
    .X(net3325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2937 (.A(\line_cache[314][2] ),
    .X(net3326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2938 (.A(\line_cache[156][3] ),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2939 (.A(\line_cache[300][2] ),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_04798_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2940 (.A(\line_cache[294][4] ),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2941 (.A(\line_cache[129][4] ),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2942 (.A(\line_cache[18][2] ),
    .X(net3331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2943 (.A(\line_cache[291][3] ),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2944 (.A(\line_cache[115][6] ),
    .X(net3333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2945 (.A(\line_cache[52][3] ),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2946 (.A(\line_cache[301][7] ),
    .X(net3335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2947 (.A(\line_cache[198][0] ),
    .X(net3336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2948 (.A(\line_cache[146][3] ),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2949 (.A(\line_cache[286][1] ),
    .X(net3338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\line_cache[167][1] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2950 (.A(\line_cache[54][4] ),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2951 (.A(\line_cache[282][4] ),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2952 (.A(\line_cache[219][2] ),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2953 (.A(\line_cache[294][2] ),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2954 (.A(\line_cache[57][0] ),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2955 (.A(\line_cache[84][1] ),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2956 (.A(\line_cache[66][4] ),
    .X(net3345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2957 (.A(\line_cache[118][7] ),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2958 (.A(\line_cache[72][6] ),
    .X(net3347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2959 (.A(\line_cache[248][2] ),
    .X(net3348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_06079_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2960 (.A(\line_cache[286][4] ),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2961 (.A(\line_cache[202][1] ),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2962 (.A(\line_cache[52][1] ),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2963 (.A(\line_cache[264][6] ),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2964 (.A(\line_cache[293][5] ),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2965 (.A(\line_cache[298][1] ),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2966 (.A(\line_cache[55][7] ),
    .X(net3355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2967 (.A(\line_cache[248][1] ),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2968 (.A(\line_cache[64][5] ),
    .X(net3357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2969 (.A(\line_cache[218][0] ),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\line_cache[267][0] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2970 (.A(\line_cache[113][0] ),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2971 (.A(\line_cache[57][7] ),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2972 (.A(\line_cache[67][3] ),
    .X(net3361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2973 (.A(\line_cache[213][1] ),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2974 (.A(\line_cache[236][4] ),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2975 (.A(\line_cache[299][1] ),
    .X(net3364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2976 (.A(\line_cache[233][6] ),
    .X(net3365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2977 (.A(\line_cache[209][4] ),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2978 (.A(\line_cache[25][6] ),
    .X(net3367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2979 (.A(\line_cache[146][4] ),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_07911_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2980 (.A(\line_cache[197][5] ),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2981 (.A(\line_cache[84][7] ),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2982 (.A(\line_cache[58][1] ),
    .X(net3371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2983 (.A(\line_cache[311][0] ),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2984 (.A(\line_cache[16][4] ),
    .X(net3373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2985 (.A(\line_cache[144][5] ),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2986 (.A(\line_cache[229][2] ),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2987 (.A(\line_cache[83][6] ),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2988 (.A(\line_cache[218][2] ),
    .X(net3377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2989 (.A(\line_cache[82][6] ),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\line_cache[158][2] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2990 (.A(\line_cache[47][0] ),
    .X(net3379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2991 (.A(\line_cache[254][1] ),
    .X(net3380));
 sky130_fd_sc_hd__buf_1 hold2992 (.A(\line_cache_idx[5] ),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2993 (.A(_00031_),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2994 (.A(\line_cache[129][3] ),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2995 (.A(\line_cache[305][2] ),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2996 (.A(\line_cache[298][4] ),
    .X(net3385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2997 (.A(\line_cache[197][6] ),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2998 (.A(\line_cache[276][3] ),
    .X(net3387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2999 (.A(\line_cache[131][3] ),
    .X(net3388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\line_cache[223][1] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_04868_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_05918_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3000 (.A(\line_cache[20][1] ),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3001 (.A(\line_cache[232][2] ),
    .X(net3390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3002 (.A(\line_cache[59][2] ),
    .X(net3391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3003 (.A(\line_cache[308][1] ),
    .X(net3392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3004 (.A(\line_cache[160][5] ),
    .X(net3393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3005 (.A(\line_cache[67][2] ),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3006 (.A(\line_cache[210][2] ),
    .X(net3395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3007 (.A(\line_cache[68][1] ),
    .X(net3396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3008 (.A(\line_cache[248][5] ),
    .X(net3397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3009 (.A(\line_cache[147][5] ),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\line_cache[262][4] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3010 (.A(\line_cache[67][4] ),
    .X(net3399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3011 (.A(\line_cache[20][5] ),
    .X(net3400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3012 (.A(\line_cache[203][3] ),
    .X(net3401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3013 (.A(\line_cache[114][1] ),
    .X(net3402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3014 (.A(\line_cache[62][0] ),
    .X(net3403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3015 (.A(\line_cache[84][5] ),
    .X(net3404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3016 (.A(\line_cache[116][5] ),
    .X(net3405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3017 (.A(\line_cache[76][4] ),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3018 (.A(\line_cache[38][6] ),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3019 (.A(\line_cache[233][5] ),
    .X(net3408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_07829_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3020 (.A(\line_cache[35][0] ),
    .X(net3409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3021 (.A(\line_cache[283][2] ),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3022 (.A(\line_cache[47][5] ),
    .X(net3411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3023 (.A(\line_cache[23][7] ),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3024 (.A(\line_cache[277][0] ),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3025 (.A(\line_cache[219][6] ),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3026 (.A(\line_cache[64][2] ),
    .X(net3415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3027 (.A(\line_cache[316][3] ),
    .X(net3416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3028 (.A(\line_cache[230][0] ),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3029 (.A(\line_cache[112][3] ),
    .X(net3418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\line_cache[139][0] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3030 (.A(\line_cache[208][1] ),
    .X(net3419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3031 (.A(\line_cache[46][1] ),
    .X(net3420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3032 (.A(\line_cache[68][4] ),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3033 (.A(\line_cache[160][6] ),
    .X(net3422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3034 (.A(\line_cache[214][1] ),
    .X(net3423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3035 (.A(\line_cache[136][5] ),
    .X(net3424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(\line_cache[268][0] ),
    .X(net3425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3037 (.A(\line_cache[318][7] ),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3038 (.A(\line_cache[277][7] ),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3039 (.A(\line_cache[172][2] ),
    .X(net3428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_05547_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3040 (.A(\line_cache[309][3] ),
    .X(net3429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3041 (.A(\line_cache[120][4] ),
    .X(net3430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3042 (.A(\line_cache[290][6] ),
    .X(net3431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3043 (.A(\line_cache[219][3] ),
    .X(net3432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3044 (.A(\line_cache[140][5] ),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3045 (.A(\line_cache[0][4] ),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3046 (.A(\line_cache[274][4] ),
    .X(net3435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3047 (.A(\line_cache[112][6] ),
    .X(net3436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3048 (.A(\line_cache[47][3] ),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3049 (.A(\line_cache[130][5] ),
    .X(net3438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\line_cache[125][4] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3050 (.A(\line_cache[224][2] ),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3051 (.A(\line_cache[217][6] ),
    .X(net3440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3052 (.A(\line_cache[33][4] ),
    .X(net3441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3053 (.A(\line_cache[72][2] ),
    .X(net3442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3054 (.A(\line_cache[172][0] ),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3055 (.A(\line_cache[20][0] ),
    .X(net3444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3056 (.A(\line_cache[200][0] ),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3057 (.A(\line_cache[61][4] ),
    .X(net3446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3058 (.A(\line_cache[231][1] ),
    .X(net3447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3059 (.A(\line_cache[176][0] ),
    .X(net3448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_05274_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3060 (.A(\line_cache[283][6] ),
    .X(net3449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3061 (.A(\line_cache[122][4] ),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3062 (.A(\res_v_counter[6] ),
    .X(net3451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3063 (.A(_00167_),
    .X(net3452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3064 (.A(\line_cache[32][0] ),
    .X(net3453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3065 (.A(\line_cache[290][0] ),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3066 (.A(\line_cache[285][6] ),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3067 (.A(\line_cache[67][5] ),
    .X(net3456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3068 (.A(\line_cache[318][2] ),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3069 (.A(\line_cache[219][0] ),
    .X(net3458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\line_cache[262][3] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3070 (.A(\line_cache[214][2] ),
    .X(net3459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3071 (.A(\line_cache[260][7] ),
    .X(net3460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3072 (.A(\line_cache[162][1] ),
    .X(net3461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3073 (.A(\line_cache[112][5] ),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3074 (.A(\line_cache[27][5] ),
    .X(net3463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3075 (.A(\line_cache[121][2] ),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3076 (.A(\line_cache[116][0] ),
    .X(net3465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3077 (.A(\line_cache[293][2] ),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3078 (.A(\line_cache[83][0] ),
    .X(net3467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3079 (.A(\line_cache[312][6] ),
    .X(net3468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_07827_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3080 (.A(\line_cache[17][0] ),
    .X(net3469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3081 (.A(\line_cache[115][0] ),
    .X(net3470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3082 (.A(\line_cache[100][2] ),
    .X(net3471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3083 (.A(\line_cache[98][1] ),
    .X(net3472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3084 (.A(\line_cache[234][1] ),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3085 (.A(\line_cache[277][1] ),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3086 (.A(\line_cache[34][1] ),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3087 (.A(\line_cache[27][7] ),
    .X(net3476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3088 (.A(\line_cache[282][0] ),
    .X(net3477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3089 (.A(\line_cache[300][6] ),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\line_cache[90][7] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3090 (.A(\line_cache[312][1] ),
    .X(net3479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3091 (.A(\line_cache[57][2] ),
    .X(net3480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3092 (.A(\line_cache[23][4] ),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3093 (.A(\line_cache[195][1] ),
    .X(net3482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3094 (.A(\line_cache[272][7] ),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3095 (.A(\line_cache[315][1] ),
    .X(net3484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3096 (.A(\line_cache[274][1] ),
    .X(net3485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3097 (.A(\base_v_sync[0] ),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3098 (.A(\line_cache[28][4] ),
    .X(net3487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3099 (.A(\line_cache[80][5] ),
    .X(net3488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\line_cache[243][5] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_04611_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3100 (.A(\line_cache[136][4] ),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3101 (.A(\line_cache[296][7] ),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3102 (.A(\line_cache[83][2] ),
    .X(net3491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3103 (.A(\line_cache[68][2] ),
    .X(net3492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3104 (.A(\line_cache[209][5] ),
    .X(net3493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3105 (.A(net106),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3106 (.A(_00049_),
    .X(net3495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3107 (.A(\line_cache[275][1] ),
    .X(net3496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3108 (.A(net104),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3109 (.A(_00047_),
    .X(net3498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\line_cache[89][3] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3110 (.A(\line_cache[124][7] ),
    .X(net3499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3111 (.A(\line_cache[22][3] ),
    .X(net3500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3112 (.A(\line_cache[17][3] ),
    .X(net3501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3113 (.A(\line_cache[118][2] ),
    .X(net3502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3114 (.A(\line_cache[113][3] ),
    .X(net3503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3115 (.A(\line_cache[197][4] ),
    .X(net3504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3116 (.A(\line_cache[55][1] ),
    .X(net3505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3117 (.A(\line_cache[318][6] ),
    .X(net3506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3118 (.A(\line_cache[253][1] ),
    .X(net3507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3119 (.A(\line_cache[114][5] ),
    .X(net3508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_04580_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3120 (.A(\line_cache[188][5] ),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3121 (.A(\line_cache[115][7] ),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3122 (.A(\line_cache[198][6] ),
    .X(net3511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3123 (.A(\line_cache[17][4] ),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3124 (.A(\line_cache[184][5] ),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3125 (.A(\line_cache[80][3] ),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3126 (.A(\line_cache[45][6] ),
    .X(net3515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3127 (.A(\line_cache[196][5] ),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3128 (.A(\line_cache[122][6] ),
    .X(net3517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3129 (.A(\line_cache[268][7] ),
    .X(net3518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\line_cache[158][5] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3130 (.A(\line_cache[47][2] ),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3131 (.A(\line_cache[117][2] ),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3132 (.A(\line_cache[304][5] ),
    .X(net3521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3133 (.A(\line_cache[130][2] ),
    .X(net3522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3134 (.A(\line_cache[30][7] ),
    .X(net3523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3135 (.A(\line_cache[44][4] ),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3136 (.A(\line_cache[50][3] ),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3137 (.A(\line_cache[88][3] ),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3138 (.A(\line_cache[232][7] ),
    .X(net3527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3139 (.A(\line_cache[119][2] ),
    .X(net3528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_05924_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3140 (.A(\line_cache[277][6] ),
    .X(net3529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3141 (.A(\line_cache[312][0] ),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3142 (.A(\line_cache[318][5] ),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3143 (.A(\line_cache[92][2] ),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3144 (.A(\line_cache[304][2] ),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3145 (.A(\line_cache[290][3] ),
    .X(net3534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3146 (.A(\line_cache[254][4] ),
    .X(net3535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3147 (.A(\line_cache[248][6] ),
    .X(net3536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3148 (.A(\line_cache[58][2] ),
    .X(net3537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3149 (.A(\line_cache[219][1] ),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\line_cache[262][1] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3150 (.A(\line_cache[202][6] ),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3151 (.A(\line_cache[318][4] ),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3152 (.A(\line_cache[272][3] ),
    .X(net3541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3153 (.A(\line_cache[295][4] ),
    .X(net3542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3154 (.A(\line_cache[122][7] ),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3155 (.A(\line_cache[31][4] ),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3156 (.A(\line_cache[136][1] ),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3157 (.A(\line_cache[295][3] ),
    .X(net3546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3158 (.A(\line_cache[268][5] ),
    .X(net3547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3159 (.A(\line_cache[235][1] ),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_07823_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3160 (.A(\line_cache[120][0] ),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3161 (.A(\line_cache[44][5] ),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3162 (.A(\line_cache[202][4] ),
    .X(net3551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3163 (.A(\line_cache[199][4] ),
    .X(net3552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3164 (.A(\line_cache[295][5] ),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3165 (.A(\line_cache[188][4] ),
    .X(net3554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3166 (.A(\line_cache[72][0] ),
    .X(net3555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3167 (.A(\line_cache[98][6] ),
    .X(net3556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3168 (.A(net95),
    .X(net3557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3169 (.A(_00038_),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\line_cache[191][4] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3170 (.A(\line_cache[164][0] ),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3171 (.A(\line_cache[199][5] ),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3172 (.A(\line_cache[274][3] ),
    .X(net3561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3173 (.A(\line_cache[118][6] ),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3174 (.A(\line_cache[234][7] ),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3175 (.A(\line_cache[198][2] ),
    .X(net3564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3176 (.A(\line_cache[39][1] ),
    .X(net3565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3177 (.A(\line_cache[147][1] ),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3178 (.A(\line_cache[230][2] ),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3179 (.A(\line_cache[264][4] ),
    .X(net3568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_06523_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3180 (.A(\line_cache[83][7] ),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3181 (.A(\line_cache[281][3] ),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3182 (.A(\line_cache[292][3] ),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3183 (.A(\line_cache[17][1] ),
    .X(net3572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3184 (.A(\line_cache[128][5] ),
    .X(net3573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3185 (.A(\line_cache[210][4] ),
    .X(net3574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3186 (.A(\line_cache[194][1] ),
    .X(net3575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3187 (.A(\line_cache[309][2] ),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3188 (.A(\line_cache[82][4] ),
    .X(net3577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3189 (.A(\line_cache[131][1] ),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\line_cache[155][0] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3190 (.A(\line_cache[204][4] ),
    .X(net3579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3191 (.A(\line_cache[16][0] ),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3192 (.A(\line_cache[62][5] ),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3193 (.A(\line_cache[57][6] ),
    .X(net3582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3194 (.A(\line_cache[172][6] ),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3195 (.A(\line_cache[188][1] ),
    .X(net3584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3196 (.A(\line_cache[213][2] ),
    .X(net3585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3197 (.A(\line_cache[253][6] ),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3198 (.A(\line_cache[183][6] ),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3199 (.A(\line_cache[57][1] ),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_07477_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_05856_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3200 (.A(\line_cache[198][4] ),
    .X(net3589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3201 (.A(\line_cache[218][5] ),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3202 (.A(\line_cache[162][0] ),
    .X(net3591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3203 (.A(\line_cache[204][7] ),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3204 (.A(\line_cache[148][2] ),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3205 (.A(\line_cache[217][7] ),
    .X(net3594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3206 (.A(\base_v_fporch[0] ),
    .X(net3595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3207 (.A(\line_cache[122][3] ),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3208 (.A(\line_cache[156][5] ),
    .X(net3597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3209 (.A(\line_cache[215][6] ),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\line_cache[138][3] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3210 (.A(\line_cache[199][1] ),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3211 (.A(\line_cache[318][1] ),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3212 (.A(\line_cache[61][5] ),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3213 (.A(\line_cache[183][7] ),
    .X(net3602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3214 (.A(\line_cache[25][3] ),
    .X(net3603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3215 (.A(\line_cache[48][7] ),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3216 (.A(\line_cache[252][5] ),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3217 (.A(\line_cache[163][2] ),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3218 (.A(net116),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3219 (.A(_00059_),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_05532_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3220 (.A(\line_cache[304][1] ),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3221 (.A(\line_cache[96][2] ),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3222 (.A(\line_cache[203][4] ),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3223 (.A(\line_cache[162][6] ),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3224 (.A(\line_cache[72][4] ),
    .X(net3613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3225 (.A(\line_cache[317][7] ),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3226 (.A(\line_cache[152][0] ),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3227 (.A(\line_cache[183][3] ),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3228 (.A(\line_cache[44][7] ),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3229 (.A(net101),
    .X(net3618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\line_cache[137][3] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3230 (.A(_00044_),
    .X(net3619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3231 (.A(\line_cache[264][2] ),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3232 (.A(\line_cache[98][2] ),
    .X(net3621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3233 (.A(\line_cache[83][4] ),
    .X(net3622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3234 (.A(\line_cache[319][4] ),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3235 (.A(net99),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3236 (.A(_00042_),
    .X(net3625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3237 (.A(\line_cache[186][6] ),
    .X(net3626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3238 (.A(\line_cache[108][1] ),
    .X(net3627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3239 (.A(\line_cache[164][1] ),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_05503_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3240 (.A(\line_cache[215][3] ),
    .X(net3629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3241 (.A(\line_cache[61][7] ),
    .X(net3630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3242 (.A(\line_cache[230][4] ),
    .X(net3631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3243 (.A(\line_cache[285][1] ),
    .X(net3632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3244 (.A(\line_cache[179][4] ),
    .X(net3633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3245 (.A(\line_cache[230][3] ),
    .X(net3634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3246 (.A(\line_cache[178][1] ),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3247 (.A(\line_cache[44][0] ),
    .X(net3636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3248 (.A(\line_cache[144][6] ),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3249 (.A(\res_h_counter[3] ),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\line_cache[267][3] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3250 (.A(_00154_),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3251 (.A(\line_cache[163][0] ),
    .X(net3640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3252 (.A(\line_cache[234][0] ),
    .X(net3641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3253 (.A(\line_cache[186][7] ),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3254 (.A(\line_cache[319][2] ),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3255 (.A(\line_cache[145][2] ),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3256 (.A(\line_cache[132][6] ),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3257 (.A(\line_cache[145][6] ),
    .X(net3646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3258 (.A(\line_cache[253][4] ),
    .X(net3647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3259 (.A(\line_cache[219][7] ),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_07917_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3260 (.A(\line_cache[132][2] ),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3261 (.A(\line_cache[58][3] ),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3262 (.A(\line_cache[202][5] ),
    .X(net3651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3263 (.A(\line_cache[25][4] ),
    .X(net3652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3264 (.A(\line_cache[235][7] ),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3265 (.A(\line_cache[92][5] ),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3266 (.A(\line_cache[305][6] ),
    .X(net3655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3267 (.A(\line_cache[176][2] ),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3268 (.A(\line_cache[183][5] ),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3269 (.A(\line_cache[44][6] ),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\line_cache[271][4] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3270 (.A(\line_cache[253][3] ),
    .X(net3659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3271 (.A(net108),
    .X(net3660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3272 (.A(_00051_),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3273 (.A(\line_cache[281][6] ),
    .X(net3662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3274 (.A(\line_cache[179][6] ),
    .X(net3663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3275 (.A(\line_cache[286][3] ),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3276 (.A(\line_cache[268][6] ),
    .X(net3665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3277 (.A(\line_cache[208][0] ),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3278 (.A(\line_cache[318][0] ),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3279 (.A(\line_cache[39][3] ),
    .X(net3668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_07991_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3280 (.A(\line_cache[24][3] ),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3281 (.A(\line_cache[187][6] ),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3282 (.A(\line_cache[255][3] ),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3283 (.A(\line_cache[179][2] ),
    .X(net3672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3284 (.A(\line_cache[255][1] ),
    .X(net3673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3285 (.A(\line_cache[183][2] ),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3286 (.A(\line_cache[83][5] ),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3287 (.A(\line_cache[43][5] ),
    .X(net3676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3288 (.A(\line_cache[156][7] ),
    .X(net3677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3289 (.A(\line_cache[113][4] ),
    .X(net3678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\line_cache[93][3] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3290 (.A(\line_cache[47][7] ),
    .X(net3679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3291 (.A(\line_cache[39][0] ),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3292 (.A(\line_cache[40][0] ),
    .X(net3681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3293 (.A(\line_cache[164][6] ),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3294 (.A(\line_cache[43][4] ),
    .X(net3683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3295 (.A(\line_cache[98][4] ),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3296 (.A(\line_cache[319][3] ),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3297 (.A(\line_cache[178][6] ),
    .X(net3686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3298 (.A(\line_cache[203][6] ),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3299 (.A(\line_cache[25][1] ),
    .X(net3688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\line_cache[267][5] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_04655_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3300 (.A(\line_cache[47][4] ),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3301 (.A(\line_cache[280][5] ),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3302 (.A(\line_cache[285][7] ),
    .X(net3691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3303 (.A(\line_cache[319][7] ),
    .X(net3692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3304 (.A(\line_cache[254][6] ),
    .X(net3693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3305 (.A(\line_cache[40][3] ),
    .X(net3694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3306 (.A(\line_cache[119][7] ),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3307 (.A(\line_cache[39][7] ),
    .X(net3696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3308 (.A(\line_cache[16][5] ),
    .X(net3697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3309 (.A(\base_h_fporch[0] ),
    .X(net3698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\line_cache[94][2] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3310 (.A(\line_cache[253][2] ),
    .X(net3699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3311 (.A(\line_cache[59][1] ),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3312 (.A(\base_h_sync[0] ),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3313 (.A(\line_cache[187][7] ),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3314 (.A(\line_cache[24][1] ),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3315 (.A(\res_v_active[5] ),
    .X(net3704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3316 (.A(\line_cache[40][1] ),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3317 (.A(\line_cache[148][0] ),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3318 (.A(\base_h_fporch[4] ),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3319 (.A(\line_cache[235][3] ),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_04674_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3320 (.A(\line_cache[286][5] ),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3321 (.A(\line_cache[172][7] ),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3322 (.A(\line_cache[317][1] ),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3323 (.A(\line_cache[39][4] ),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3324 (.A(\base_v_counter[9] ),
    .X(net3713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3325 (.A(_12959_),
    .X(net3714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3326 (.A(_00150_),
    .X(net3715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3327 (.A(\line_cache[144][2] ),
    .X(net3716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3328 (.A(\line_cache[162][2] ),
    .X(net3717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3329 (.A(\line_cache[152][2] ),
    .X(net3718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\line_cache[175][1] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3330 (.A(\line_cache[168][0] ),
    .X(net3719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3331 (.A(\line_cache[235][2] ),
    .X(net3720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3332 (.A(\line_cache[202][0] ),
    .X(net3721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3333 (.A(\line_cache[178][5] ),
    .X(net3722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3334 (.A(\line_cache[179][1] ),
    .X(net3723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3335 (.A(\line_cache[210][0] ),
    .X(net3724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3336 (.A(\line_cache[204][3] ),
    .X(net3725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3337 (.A(\line_cache[184][1] ),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3338 (.A(\line_cache[210][1] ),
    .X(net3727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3339 (.A(\line_cache[43][6] ),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_06226_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3340 (.A(\line_cache[120][7] ),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3341 (.A(\line_cache[92][3] ),
    .X(net3730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3342 (.A(\line_cache[281][1] ),
    .X(net3731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3343 (.A(\line_cache[24][4] ),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3344 (.A(\line_cache[179][5] ),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3345 (.A(\line_cache[209][0] ),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3346 (.A(\resolution[1] ),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3347 (.A(\line_cache[43][7] ),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3348 (.A(\line_cache[220][2] ),
    .X(net3737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3349 (.A(\resolution[3] ),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\line_cache[75][7] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3350 (.A(\line_cache[215][1] ),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3351 (.A(\line_cache[281][5] ),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3352 (.A(\line_cache[40][4] ),
    .X(net3741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3353 (.A(\line_cache[43][0] ),
    .X(net3742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3354 (.A(\line_cache[178][2] ),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3355 (.A(\line_cache[215][5] ),
    .X(net3744));
 sky130_fd_sc_hd__buf_1 hold3356 (.A(\res_h_counter[2] ),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3357 (.A(_00153_),
    .X(net3746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3358 (.A(\res_v_active[4] ),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3359 (.A(\line_cache[254][5] ),
    .X(net3748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_04331_),
    .X(net725));
 sky130_fd_sc_hd__buf_1 hold3360 (.A(\res_v_counter[3] ),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3361 (.A(_00164_),
    .X(net3750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3362 (.A(\line_cache[235][6] ),
    .X(net3751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3363 (.A(\line_cache[43][3] ),
    .X(net3752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3364 (.A(\line_cache[44][3] ),
    .X(net3753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3365 (.A(\line_cache[178][4] ),
    .X(net3754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3366 (.A(\line_cache[218][6] ),
    .X(net3755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3367 (.A(\prescaler[2] ),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3368 (.A(\line_cache[319][0] ),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3369 (.A(\res_v_active[2] ),
    .X(net3758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\line_cache[137][0] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3370 (.A(\line_cache[215][4] ),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3371 (.A(\line_cache[99][4] ),
    .X(net3760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3372 (.A(\line_cache[305][7] ),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3373 (.A(\line_cache[319][5] ),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3374 (.A(\resolution[2] ),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3375 (.A(net96),
    .X(net3764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3376 (.A(_00039_),
    .X(net3765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3377 (.A(\line_cache[253][5] ),
    .X(net3766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3378 (.A(\line_cache[40][7] ),
    .X(net3767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3379 (.A(net102),
    .X(net3768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_05490_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3380 (.A(_00045_),
    .X(net3769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3381 (.A(\line_cache[184][6] ),
    .X(net3770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3382 (.A(\line_cache[319][6] ),
    .X(net3771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3383 (.A(\line_cache[43][1] ),
    .X(net3772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3384 (.A(\res_h_counter[0] ),
    .X(net3773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3385 (.A(_00151_),
    .X(net3774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3386 (.A(\line_cache[286][6] ),
    .X(net3775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3387 (.A(\line_cache[305][0] ),
    .X(net3776));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3388 (.A(\res_v_counter[5] ),
    .X(net3777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3389 (.A(_00166_),
    .X(net3778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\line_cache[103][4] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3390 (.A(\line_cache[255][4] ),
    .X(net3779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3391 (.A(\res_v_active[3] ),
    .X(net3780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3392 (.A(\line_cache[61][6] ),
    .X(net3781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3393 (.A(\line_cache[44][1] ),
    .X(net3782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3394 (.A(\line_cache[97][4] ),
    .X(net3783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3395 (.A(\base_v_counter[3] ),
    .X(net3784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3396 (.A(_12895_),
    .X(net3785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3397 (.A(_00144_),
    .X(net3786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3398 (.A(\line_cache[235][4] ),
    .X(net3787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3399 (.A(\line_cache[264][1] ),
    .X(net3788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_07921_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_04841_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3400 (.A(\line_cache[200][2] ),
    .X(net3789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3401 (.A(net105),
    .X(net3790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3402 (.A(_00048_),
    .X(net3791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3403 (.A(net107),
    .X(net3792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3404 (.A(_00050_),
    .X(net3793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3405 (.A(\line_cache[254][3] ),
    .X(net3794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3406 (.A(\line_cache[235][5] ),
    .X(net3795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3407 (.A(\line_cache[116][7] ),
    .X(net3796));
 sky130_fd_sc_hd__clkbuf_2 hold3408 (.A(\base_v_counter[4] ),
    .X(net3797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3409 (.A(_12907_),
    .X(net3798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\line_cache[11][7] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3410 (.A(_00145_),
    .X(net3799));
 sky130_fd_sc_hd__buf_1 hold3411 (.A(\base_v_counter[1] ),
    .X(net3800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3412 (.A(_12856_),
    .X(net3801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3413 (.A(_00142_),
    .X(net3802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3414 (.A(\line_cache[215][2] ),
    .X(net3803));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3415 (.A(\res_v_counter[2] ),
    .X(net3804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3416 (.A(_00163_),
    .X(net3805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3417 (.A(\line_cache[116][6] ),
    .X(net3806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3418 (.A(\line_cache[255][2] ),
    .X(net3807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3419 (.A(\line_cache[31][6] ),
    .X(net3808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_03131_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3420 (.A(\line_cache[172][3] ),
    .X(net3809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3421 (.A(\line_cache[319][1] ),
    .X(net3810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3422 (.A(\line_cache[108][3] ),
    .X(net3811));
 sky130_fd_sc_hd__buf_1 hold3423 (.A(\base_v_counter[6] ),
    .X(net3812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3424 (.A(_12930_),
    .X(net3813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3425 (.A(_00147_),
    .X(net3814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3426 (.A(\base_v_active[8] ),
    .X(net3815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3427 (.A(\base_h_bporch[0] ),
    .X(net3816));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3428 (.A(\base_v_counter[5] ),
    .X(net3817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3429 (.A(_12918_),
    .X(net3818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\line_cache[189][4] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3430 (.A(_00146_),
    .X(net3819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3431 (.A(\res_v_active[6] ),
    .X(net3820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3432 (.A(net103),
    .X(net3821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3433 (.A(_00046_),
    .X(net3822));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3434 (.A(\base_v_counter[8] ),
    .X(net3823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3435 (.A(_12952_),
    .X(net3824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3436 (.A(\line_cache[31][1] ),
    .X(net3825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3437 (.A(\line_cache[203][1] ),
    .X(net3826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3438 (.A(\line_cache[204][1] ),
    .X(net3827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3439 (.A(\line_cache[204][5] ),
    .X(net3828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_06486_),
    .X(net733));
 sky130_fd_sc_hd__buf_1 hold3440 (.A(\res_v_counter[0] ),
    .X(net3829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3441 (.A(_00161_),
    .X(net3830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3442 (.A(\line_cache[286][0] ),
    .X(net3831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3443 (.A(\base_h_fporch[2] ),
    .X(net3832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3444 (.A(\line_cache[31][2] ),
    .X(net3833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3445 (.A(\base_h_sync[4] ),
    .X(net3834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3446 (.A(\base_v_active[1] ),
    .X(net3835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3447 (.A(\res_v_counter[7] ),
    .X(net3836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3448 (.A(_00168_),
    .X(net3837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3449 (.A(\base_v_fporch[2] ),
    .X(net3838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\line_cache[89][1] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3450 (.A(\line_cache[120][6] ),
    .X(net3839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3451 (.A(\line_cache[203][0] ),
    .X(net3840));
 sky130_fd_sc_hd__buf_1 hold3452 (.A(net113),
    .X(net3841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3453 (.A(_12403_),
    .X(net3842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3454 (.A(_00056_),
    .X(net3843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3455 (.A(\base_h_active[7] ),
    .X(net3844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3456 (.A(\line_cache[31][3] ),
    .X(net3845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3457 (.A(net109),
    .X(net3846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3458 (.A(_12384_),
    .X(net3847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3459 (.A(_00052_),
    .X(net3848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_04574_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3460 (.A(\line_cache[31][5] ),
    .X(net3849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3461 (.A(\base_v_active[2] ),
    .X(net3850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3462 (.A(\line_cache[31][0] ),
    .X(net3851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3463 (.A(\base_v_fporch[1] ),
    .X(net3852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3464 (.A(\res_v_active[1] ),
    .X(net3853));
 sky130_fd_sc_hd__buf_1 hold3465 (.A(net97),
    .X(net3854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3466 (.A(_12349_),
    .X(net3855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3467 (.A(_00040_),
    .X(net3856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3468 (.A(\base_h_sync[5] ),
    .X(net3857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3469 (.A(\line_cache[286][2] ),
    .X(net3858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\line_cache[69][5] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3470 (.A(\line_cache[286][7] ),
    .X(net3859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3471 (.A(net115),
    .X(net3860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3472 (.A(_12409_),
    .X(net3861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3473 (.A(_00058_),
    .X(net3862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3474 (.A(\res_v_active[7] ),
    .X(net3863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3475 (.A(\line_cache[162][4] ),
    .X(net3864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3476 (.A(\line_cache[203][5] ),
    .X(net3865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3477 (.A(\prescaler[1] ),
    .X(net3866));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3478 (.A(\res_h_counter[1] ),
    .X(net3867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3479 (.A(_00152_),
    .X(net3868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_04216_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3480 (.A(\line_cache[186][0] ),
    .X(net3869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3481 (.A(\base_h_active[9] ),
    .X(net3870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3482 (.A(\line_cache[44][2] ),
    .X(net3871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3483 (.A(\prescaler_counter[6] ),
    .X(net3872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3484 (.A(_09521_),
    .X(net3873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3485 (.A(_09522_),
    .X(net3874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3486 (.A(\line_cache[39][5] ),
    .X(net3875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3487 (.A(\base_v_sync[1] ),
    .X(net3876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3488 (.A(\base_h_fporch[1] ),
    .X(net3877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3489 (.A(\line_cache[39][6] ),
    .X(net3878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\line_cache[263][1] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3490 (.A(\line_cache[163][4] ),
    .X(net3879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3491 (.A(\res_v_active[0] ),
    .X(net3880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3492 (.A(\base_h_bporch[3] ),
    .X(net3881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3493 (.A(\line_cache[40][6] ),
    .X(net3882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3494 (.A(\line_cache[287][3] ),
    .X(net3883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3495 (.A(\base_h_bporch[5] ),
    .X(net3884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3496 (.A(net125),
    .X(net3885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3497 (.A(_08826_),
    .X(net3886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3498 (.A(\base_h_fporch[3] ),
    .X(net3887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3499 (.A(\prescaler_counter[5] ),
    .X(net3888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\line_cache[1][1] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_07839_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3500 (.A(_09517_),
    .X(net3889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3501 (.A(_09518_),
    .X(net3890));
 sky130_fd_sc_hd__buf_1 hold3502 (.A(\prescaler[3] ),
    .X(net3891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3503 (.A(\line_cache[43][2] ),
    .X(net3892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3504 (.A(\base_h_sync[3] ),
    .X(net3893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3505 (.A(\base_h_bporch[4] ),
    .X(net3894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3506 (.A(\base_h_active[2] ),
    .X(net3895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3507 (.A(\base_h_active[4] ),
    .X(net3896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3508 (.A(\base_v_bporch[3] ),
    .X(net3897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3509 (.A(\line_cache[187][0] ),
    .X(net3898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\line_cache[238][6] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3510 (.A(\line_cache[31][7] ),
    .X(net3899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3511 (.A(net94),
    .X(net3900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3512 (.A(_00037_),
    .X(net3901));
 sky130_fd_sc_hd__buf_1 hold3513 (.A(\res_h_counter[5] ),
    .X(net3902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3514 (.A(_00156_),
    .X(net3903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3515 (.A(\base_v_bporch[1] ),
    .X(net3904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3516 (.A(\base_v_sync[2] ),
    .X(net3905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3517 (.A(\base_v_active[7] ),
    .X(net3906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3518 (.A(\resolution[0] ),
    .X(net3907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3519 (.A(\base_v_active[5] ),
    .X(net3908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_07389_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3520 (.A(\line_cache[287][5] ),
    .X(net3909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3521 (.A(\res_h_active[1] ),
    .X(net3910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3522 (.A(\base_h_active[8] ),
    .X(net3911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3523 (.A(\line_cache[40][5] ),
    .X(net3912));
 sky130_fd_sc_hd__clkbuf_2 hold3524 (.A(\line_cache_idx[7] ),
    .X(net3913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3525 (.A(_00033_),
    .X(net3914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3526 (.A(\res_h_counter[7] ),
    .X(net3915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3527 (.A(_00158_),
    .X(net3916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3528 (.A(\line_cache[287][7] ),
    .X(net3917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3529 (.A(\base_h_sync[6] ),
    .X(net3918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\line_cache[250][1] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3530 (.A(\line_cache[287][4] ),
    .X(net3919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3531 (.A(\line_cache[287][6] ),
    .X(net3920));
 sky130_fd_sc_hd__buf_4 hold3532 (.A(\line_cache_idx[3] ),
    .X(net3921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3533 (.A(_00029_),
    .X(net3922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3534 (.A(\base_h_active[0] ),
    .X(net3923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3535 (.A(\line_cache[287][2] ),
    .X(net3924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3536 (.A(\line_cache[287][1] ),
    .X(net3925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3537 (.A(\base_h_sync[2] ),
    .X(net3926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3538 (.A(\base_v_active[0] ),
    .X(net3927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3539 (.A(\base_h_active[6] ),
    .X(net3928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_07599_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3540 (.A(\res_h_active[0] ),
    .X(net3929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3541 (.A(\line_cache[287][0] ),
    .X(net3930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3542 (.A(\res_h_active[3] ),
    .X(net3931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3543 (.A(\base_h_bporch[1] ),
    .X(net3932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3544 (.A(\line_cache[255][0] ),
    .X(net3933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3545 (.A(\base_h_sync[1] ),
    .X(net3934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3546 (.A(\base_h_bporch[6] ),
    .X(net3935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3547 (.A(\base_v_counter[7] ),
    .X(net3936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3548 (.A(_12942_),
    .X(net3937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3549 (.A(\base_v_active[4] ),
    .X(net3938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\line_cache[155][2] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3550 (.A(\base_v_bporch[0] ),
    .X(net3939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3551 (.A(\base_h_active[5] ),
    .X(net3940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3552 (.A(\line_cache[255][7] ),
    .X(net3941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3553 (.A(\base_h_active[1] ),
    .X(net3942));
 sky130_fd_sc_hd__buf_1 hold3554 (.A(\res_h_counter[4] ),
    .X(net3943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3555 (.A(_00155_),
    .X(net3944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3556 (.A(\res_h_active[4] ),
    .X(net3945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3557 (.A(\line_cache[255][5] ),
    .X(net3946));
 sky130_fd_sc_hd__buf_1 hold3558 (.A(\base_h_counter[9] ),
    .X(net3947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3559 (.A(_00140_),
    .X(net3948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_05860_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3560 (.A(\base_v_active[3] ),
    .X(net3949));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3561 (.A(net117),
    .X(net3950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3562 (.A(_00060_),
    .X(net3951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3563 (.A(\prescaler[0] ),
    .X(net3952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3564 (.A(\base_h_bporch[2] ),
    .X(net3953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3565 (.A(\base_v_active[6] ),
    .X(net3954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3566 (.A(\line_cache[255][6] ),
    .X(net3955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3567 (.A(net121),
    .X(net3956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3568 (.A(_00064_),
    .X(net3957));
 sky130_fd_sc_hd__buf_1 hold3569 (.A(\prescaler_counter[1] ),
    .X(net3958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\line_cache[263][6] ),
    .X(net746));
 sky130_fd_sc_hd__buf_1 hold3570 (.A(\base_h_counter[8] ),
    .X(net3959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3571 (.A(_00139_),
    .X(net3960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3572 (.A(\base_h_active[3] ),
    .X(net3961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3573 (.A(net122),
    .X(net3962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3574 (.A(_00065_),
    .X(net3963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3575 (.A(\base_v_bporch[2] ),
    .X(net3964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3576 (.A(\base_h_counter[1] ),
    .X(net3965));
 sky130_fd_sc_hd__clkbuf_2 hold3577 (.A(\res_h_active[7] ),
    .X(net3966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3578 (.A(\res_h_active[5] ),
    .X(net3967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3579 (.A(\base_h_counter[7] ),
    .X(net3968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_07850_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3580 (.A(_00138_),
    .X(net3969));
 sky130_fd_sc_hd__buf_1 hold3581 (.A(\res_h_active[6] ),
    .X(net3970));
 sky130_fd_sc_hd__clkbuf_2 hold3582 (.A(\res_h_active[8] ),
    .X(net3971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3583 (.A(\fb_read_state[1] ),
    .X(net3972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3584 (.A(_00011_),
    .X(net3973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3585 (.A(\res_h_active[2] ),
    .X(net3974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3586 (.A(net119),
    .X(net3975));
 sky130_fd_sc_hd__buf_1 hold3587 (.A(\base_h_counter[2] ),
    .X(net3976));
 sky130_fd_sc_hd__buf_1 hold3588 (.A(\fb_read_state[2] ),
    .X(net3977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3589 (.A(_00010_),
    .X(net3978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\line_cache[91][3] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3590 (.A(\prescaler_counter[8] ),
    .X(net3979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3591 (.A(_09527_),
    .X(net3980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3592 (.A(_09529_),
    .X(net3981));
 sky130_fd_sc_hd__buf_2 hold3593 (.A(\line_cache_idx[2] ),
    .X(net3982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3594 (.A(_12291_),
    .X(net3983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3595 (.A(\prescaler_counter[4] ),
    .X(net3984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3596 (.A(_09511_),
    .X(net3985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3597 (.A(_09513_),
    .X(net3986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3598 (.A(net98),
    .X(net3987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3599 (.A(\base_h_counter[3] ),
    .X(net3988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_02866_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_04619_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3600 (.A(\line_cache_idx[9] ),
    .X(net3989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3601 (.A(\base_h_counter[6] ),
    .X(net3990));
 sky130_fd_sc_hd__buf_1 hold3602 (.A(\prescaler_counter[2] ),
    .X(net3991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3603 (.A(\base_h_counter[5] ),
    .X(net3992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3604 (.A(_00136_),
    .X(net3993));
 sky130_fd_sc_hd__buf_1 hold3605 (.A(\base_h_counter[4] ),
    .X(net3994));
 sky130_fd_sc_hd__buf_1 hold3606 (.A(\line_cache_idx[4] ),
    .X(net3995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3607 (.A(net111),
    .X(net3996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3608 (.A(\prescaler_counter[7] ),
    .X(net3997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3609 (.A(net123),
    .X(net3998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\line_cache[206][5] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3610 (.A(_08828_),
    .X(net3999));
 sky130_fd_sc_hd__buf_1 hold3611 (.A(\prescaler_counter[3] ),
    .X(net4000));
 sky130_fd_sc_hd__buf_1 hold3612 (.A(\line_cache_idx[6] ),
    .X(net4001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3613 (.A(\prescaler_counter[7] ),
    .X(net4002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3614 (.A(_08835_),
    .X(net4003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3615 (.A(\prescaler_counter[0] ),
    .X(net4004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_06808_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\line_cache[190][2] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_06502_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\line_cache[95][7] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_04701_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\line_cache[261][7] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_07818_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\line_cache[243][6] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\line_cache[106][1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_07479_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\line_cache[111][7] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_04994_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\line_cache[106][4] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_04898_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\line_cache[137][2] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_05499_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\line_cache[90][5] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_04607_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\line_cache[249][0] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_04892_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_07572_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\line_cache[93][0] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_04645_),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\line_cache[125][6] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_05280_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\line_cache[89][6] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_04589_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\line_cache[93][5] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_04661_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\line_cache[1][5] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\line_cache[243][4] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_02894_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\line_cache[10][0] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_03100_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\line_cache[139][1] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_05550_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\line_cache[69][7] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_04222_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\line_cache[207][5] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_06824_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\line_cache[105][0] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_07106_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_07475_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_04865_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\line_cache[95][5] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_04697_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\line_cache[1][2] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_02873_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\line_cache[106][2] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_04894_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\line_cache[157][5] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_05905_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\line_cache[75][4] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\line_cache[1][0] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_04325_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\line_cache[174][7] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_06222_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\line_cache[150][6] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_05778_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\line_cache[166][4] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_06069_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\line_cache[101][6] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_04810_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\line_cache[250][0] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_02859_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_07597_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\line_cache[10][3] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_03107_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\line_cache[221][0] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_07063_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\line_cache[5][5] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_03017_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\line_cache[127][7] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_05317_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\line_cache[10][5] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\line_cache[246][4] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_03111_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\line_cache[91][2] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_04617_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\line_cache[70][5] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_04236_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\line_cache[171][7] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_06165_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\line_cache[143][5] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_05646_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\line_cache[271][5] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_07532_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_07993_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\line_cache[9][3] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_03085_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\line_cache[149][7] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_05763_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\line_cache[263][4] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_07846_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\line_cache[174][1] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_06209_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\line_cache[271][2] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\line_cache[77][4] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_07987_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\line_cache[10][7] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_03115_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\line_cache[7][2] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_03047_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\line_cache[150][0] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_05766_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\line_cache[174][5] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_06218_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\line_cache[87][3] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_04363_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_04545_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\line_cache[70][7] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_04240_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\line_cache[237][1] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_07355_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\line_cache[111][3] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_04986_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\line_cache[134][4] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_05448_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\line_cache[134][5] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\line_cache[1][3] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_05450_),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\line_cache[237][5] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_07367_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\line_cache[249][6] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_07591_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\line_cache[89][0] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_04571_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\line_cache[142][7] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_05634_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\line_cache[150][7] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_02880_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_05780_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\line_cache[111][0] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_04980_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\line_cache[69][6] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_04219_),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\line_cache[87][6] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_04551_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\line_cache[137][6] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_05515_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\line_cache[263][2] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\line_cache[107][3] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_07842_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\line_cache[169][4] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_06122_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\line_cache[94][1] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_04672_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\line_cache[87][4] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_04547_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\line_cache[271][7] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_07997_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\line_cache[75][6] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\line_cache[257][3] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_04913_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_04329_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\line_cache[101][0] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_04792_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\line_cache[157][3] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_05899_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\line_cache[85][3] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_04507_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\line_cache[266][1] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_07896_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\line_cache[175][0] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\line_cache[2][5] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_06224_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\line_cache[150][2] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_05770_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\line_cache[266][7] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_07909_),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\line_cache[2][1] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_02919_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\line_cache[159][7] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_05945_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\line_cache[77][2] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_02940_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_04357_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\line_cache[262][7] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_07835_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\line_cache[14][4] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_03183_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\line_cache[158][3] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_05920_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\line_cache[74][7] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_04314_),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\line_cache[143][2] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\line_cache[243][3] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_05640_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\line_cache[170][3] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_06140_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\line_cache[137][1] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_05494_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\line_cache[142][2] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_05624_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\line_cache[265][5] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_07885_),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\line_cache[79][7] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_07473_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_04406_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\line_cache[126][3] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_05292_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\line_cache[138][5] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_05538_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\line_cache[249][1] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_07575_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\line_cache[207][6] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_06826_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\line_cache[175][2] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\line_cache[106][6] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_06228_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\line_cache[153][3] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_05824_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\line_cache[103][7] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_04847_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\line_cache[250][4] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_07605_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\line_cache[79][0] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_04392_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\line_cache[5][6] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_04902_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_03020_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\line_cache[71][2] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_04246_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\line_cache[271][1] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_07985_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\line_cache[190][3] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_06504_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\line_cache[5][0] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_03001_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\line_cache[266][2] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\line_cache[258][6] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_07899_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\line_cache[105][5] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_04881_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\line_cache[263][7] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_07852_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\line_cache[109][6] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_04957_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\line_cache[142][1] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_05621_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\line_cache[78][5] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_07760_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_04386_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\line_cache[269][6] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_07961_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\line_cache[86][4] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_04530_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\line_cache[154][3] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_05846_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\line_cache[69][0] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_04201_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\line_cache[93][7] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\line_cache[258][3] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_04667_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\line_cache[169][2] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_06116_),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\line_cache[95][1] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_04688_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\line_cache[101][4] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_04804_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\line_cache[173][7] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_06204_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\line_cache[137][5] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_07732_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_07754_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_05511_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\line_cache[109][5] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_04954_),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\line_cache[85][7] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_04519_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\line_cache[174][0] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_06207_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\line_cache[257][0] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_07723_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\line_cache[78][0] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\line_cache[107][6] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_04375_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\line_cache[158][0] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_05914_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\line_cache[257][6] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_07741_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\line_cache[237][2] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_07358_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\line_cache[126][5] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_05296_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\line_cache[85][4] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_04919_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_04510_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\line_cache[237][0] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_07352_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\line_cache[138][0] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_05523_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\line_cache[91][4] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_04621_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\line_cache[262][5] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_07831_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\line_cache[9][5] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\line_cache[2][3] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_03091_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\line_cache[5][7] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_03023_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\line_cache[165][4] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_06048_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\line_cache[138][4] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_05535_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\line_cache[7][6] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_03055_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\line_cache[173][2] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_02930_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_06189_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\line_cache[157][2] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_05896_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\line_cache[157][6] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_05908_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\line_cache[75][5] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_04327_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\line_cache[165][0] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_06036_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\line_cache[109][0] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\line_cache[259][1] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_04939_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\line_cache[7][7] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_03057_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\line_cache[87][2] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_04543_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\line_cache[191][1] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_06516_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\line_cache[265][3] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_07879_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\line_cache[270][2] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_07766_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_07971_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\line_cache[223][2] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_07109_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\line_cache[191][3] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_06521_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\line_cache[94][3] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_04676_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\line_cache[265][0] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_07870_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\line_cache[173][3] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\line_cache[259][7] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_06192_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\line_cache[169][6] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_06128_),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\line_cache[126][4] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_05294_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\line_cache[151][6] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_05795_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\line_cache[141][4] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_05604_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\line_cache[170][1] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_07778_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_06136_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\line_cache[171][6] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_06163_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\line_cache[3][7] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_02982_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\line_cache[151][5] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_05793_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\line_cache[238][4] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_07385_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\line_cache[103][2] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\line_cache[246][1] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_04837_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\line_cache[149][6] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_05760_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\line_cache[135][7] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_05470_),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\line_cache[139][3] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_05557_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\line_cache[103][1] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_04835_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\line_cache[151][0] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\line_cache[78][6] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_07525_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_05782_),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\line_cache[166][3] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_06067_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\line_cache[151][3] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_05789_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\line_cache[169][3] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_06119_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\line_cache[175][4] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_06232_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\line_cache[142][3] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\line_cache[106][7] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_05626_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\line_cache[69][4] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_04213_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\line_cache[87][0] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_04538_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\line_cache[154][4] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_05848_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\line_cache[101][3] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_04801_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\line_cache[143][0] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_04904_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_05636_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\line_cache[126][2] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_05290_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\line_cache[266][6] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_07907_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\line_cache[134][2] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_05444_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\line_cache[207][3] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_06820_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\line_cache[258][4] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\line_cache[267][4] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_07756_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\line_cache[107][5] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_04917_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\line_cache[109][3] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_04948_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\line_cache[239][5] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_07403_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\line_cache[169][1] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_06112_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\line_cache[70][6] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_07919_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_04238_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\line_cache[237][3] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_07361_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\line_cache[249][7] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_07594_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\line_cache[69][2] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_04207_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\line_cache[139][7] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_05569_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\line_cache[158][6] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\line_cache[246][3] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_05926_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\line_cache[127][6] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_05315_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\line_cache[143][1] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_05638_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\line_cache[246][5] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_07534_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\line_cache[221][5] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_07079_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\line_cache[265][7] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_07530_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_07891_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\line_cache[77][3] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_04360_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\line_cache[247][5] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_07550_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\line_cache[126][7] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_05300_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\line_cache[89][7] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_04592_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\line_cache[13][6] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\line_cache[1][6] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_03169_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\line_cache[91][1] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_04615_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\line_cache[125][2] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_05268_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\line_cache[125][1] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_05264_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\line_cache[206][2] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_06802_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\line_cache[189][2] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_02901_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_06480_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\line_cache[10][4] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_03109_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\line_cache[241][0] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_07425_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\line_cache[171][1] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_06152_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\line_cache[158][1] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_05916_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\line_cache[127][3] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\line_cache[70][3] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_05309_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\line_cache[174][4] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_06216_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\line_cache[265][6] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_07888_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\line_cache[9][1] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_03079_),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\line_cache[5][3] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_03011_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\line_cache[242][5] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_04388_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_04232_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_07460_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\line_cache[137][4] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_05507_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\line_cache[157][0] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_05888_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\line_cache[174][6] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_06220_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\line_cache[173][1] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_06186_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\line_cache[95][3] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\line_cache[2][2] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_04693_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\line_cache[153][6] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_05833_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\line_cache[3][6] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_02978_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\line_cache[189][5] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_06489_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\line_cache[70][4] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_04234_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\line_cache[101][5] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_02925_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_04807_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\line_cache[110][0] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_04963_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\line_cache[79][4] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_04400_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\line_cache[165][7] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_06057_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\line_cache[87][7] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_04553_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\line_cache[270][6] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\line_cache[133][7] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_07979_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\line_cache[265][4] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_07882_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\line_cache[85][1] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_04500_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\line_cache[155][3] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_05862_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\line_cache[74][0] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_04300_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\line_cache[126][0] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_05436_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_05286_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\line_cache[143][6] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_05648_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\line_cache[245][5] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_07514_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\line_cache[127][2] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_05307_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\line_cache[110][4] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_04972_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\line_cache[101][7] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\line_cache[78][1] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_04813_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\line_cache[103][6] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_04845_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\line_cache[143][3] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_05642_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\line_cache[205][4] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_06785_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\line_cache[155][6] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_05868_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\line_cache[151][1] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_04377_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_05784_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\line_cache[135][4] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_05464_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\line_cache[110][2] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_04968_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\line_cache[5][1] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_03004_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\line_cache[247][0] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_07540_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\line_cache[250][5] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\line_cache[245][3] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_07607_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\line_cache[141][0] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_05588_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\line_cache[266][5] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_07905_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\line_cache[9][4] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_03088_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\line_cache[261][6] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_07815_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\line_cache[135][6] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_07508_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_05468_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\line_cache[150][1] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_05768_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\line_cache[79][5] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_04402_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\line_cache[206][4] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_06806_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\line_cache[242][3] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_07456_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\line_cache[90][3] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\line_cache[241][4] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_04603_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\line_cache[135][3] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_05462_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\line_cache[110][7] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_04978_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\line_cache[111][2] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_04984_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\line_cache[71][0] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_04242_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\line_cache[102][3] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\line_cache[2][6] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_07438_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_04823_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\line_cache[134][3] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_05446_),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\line_cache[13][4] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_03163_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\line_cache[125][0] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_05261_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\line_cache[191][7] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_06529_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\line_cache[269][0] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\line_cache[73][2] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_07942_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\line_cache[94][7] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_04684_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\line_cache[142][6] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_05632_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\line_cache[15][6] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_03204_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\line_cache[263][5] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_07848_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\line_cache[258][2] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_04282_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_07752_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\line_cache[86][3] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_04528_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\line_cache[173][5] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_06198_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\line_cache[257][1] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_07726_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\line_cache[191][6] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_06527_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\line_cache[155][1] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\line_cache[73][5] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_05858_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\line_cache[258][0] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_07747_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\line_cache[170][7] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_06148_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\line_cache[73][7] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_04297_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\line_cache[135][1] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_05458_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\line_cache[6][1] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_04291_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_03028_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\line_cache[6][4] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_03034_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\line_cache[259][6] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_07776_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\line_cache[103][3] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_04839_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\line_cache[79][3] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_04398_),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\line_cache[127][4] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\line_cache[258][1] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_05311_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\line_cache[165][6] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_06054_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\line_cache[141][5] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_05608_),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\line_cache[90][2] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_04601_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\line_cache[142][5] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_05630_),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\line_cache[79][2] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_07749_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_04396_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\line_cache[239][2] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_07397_),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\line_cache[3][0] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_02954_),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\line_cache[166][0] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_06060_),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\line_cache[262][6] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_07833_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\line_cache[175][3] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\line_cache[73][1] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_06230_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\line_cache[157][7] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_05911_),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\line_cache[271][0] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_07983_),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\line_cache[154][6] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_05852_),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\line_cache[167][0] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_06077_),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\line_cache[157][1] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_04278_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_05891_),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\line_cache[237][6] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_07370_),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\line_cache[103][5] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_04843_),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\line_cache[94][4] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_04678_),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\line_cache[223][3] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_07111_),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\line_cache[86][7] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\line_cache[267][7] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_04536_),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\line_cache[139][6] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_05566_),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\line_cache[110][3] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_04970_),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\line_cache[269][4] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_07955_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\line_cache[166][7] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_06075_),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\line_cache[263][0] ),
    .X(net1388));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(base_h_active_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(base_h_active_i[9]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(base_h_bporch_i[0]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(base_h_bporch_i[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(base_h_bporch_i[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(base_h_bporch_i[3]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(base_h_bporch_i[4]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(base_h_bporch_i[5]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(base_h_bporch_i[6]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(base_h_fporch_i[0]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(base_h_fporch_i[1]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(base_h_active_i[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(base_h_fporch_i[2]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(base_h_fporch_i[3]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(base_h_fporch_i[4]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(base_h_sync_i[0]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(base_h_sync_i[1]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(base_h_sync_i[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(base_h_sync_i[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(base_h_sync_i[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(base_h_sync_i[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(base_h_sync_i[6]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(base_h_active_i[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(base_v_active_i[0]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(base_v_active_i[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(base_v_active_i[2]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(base_v_active_i[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(base_v_active_i[4]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(base_v_active_i[5]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(base_v_active_i[6]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(base_v_active_i[7]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(base_v_active_i[8]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(base_v_bporch_i[0]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(base_h_active_i[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(base_v_bporch_i[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(base_v_bporch_i[2]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(base_v_bporch_i[3]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(base_v_fporch_i[0]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(base_v_fporch_i[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(base_v_fporch_i[2]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(base_v_sync_i[0]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(base_v_sync_i[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(base_v_sync_i[2]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(enable_i),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input5 (.A(base_h_active_i[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input50 (.A(mport_i[0]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(mport_i[10]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(mport_i[11]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(mport_i[12]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(mport_i[13]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(mport_i[14]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(mport_i[15]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(mport_i[16]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(mport_i[17]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(mport_i[18]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input6 (.A(base_h_active_i[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input60 (.A(mport_i[19]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(mport_i[1]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(mport_i[20]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(mport_i[21]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(mport_i[22]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(mport_i[23]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(mport_i[24]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(mport_i[25]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(mport_i[26]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(mport_i[27]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(base_h_active_i[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input70 (.A(mport_i[28]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(mport_i[29]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(mport_i[2]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(mport_i[30]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(mport_i[31]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(mport_i[33]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(mport_i[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(mport_i[4]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(mport_i[5]),
    .X(net78));
 sky130_fd_sc_hd__buf_2 input79 (.A(mport_i[6]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(base_h_active_i[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input80 (.A(mport_i[7]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(mport_i[8]),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(mport_i[9]),
    .X(net82));
 sky130_fd_sc_hd__buf_4 input83 (.A(nrst_i),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(prescaler_i[0]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(prescaler_i[1]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(prescaler_i[2]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(prescaler_i[3]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(resolution_i[0]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(resolution_i[1]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(base_h_active_i[8]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(resolution_i[2]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(resolution_i[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(mport_o[41]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(mport_o[42]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(mport_o[43]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(mport_o[44]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(mport_o[45]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(mport_o[46]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(mport_o[47]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(mport_o[48]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(mport_o[49]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(mport_o[50]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(mport_o[51]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(mport_o[52]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(mport_o[53]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(mport_o[54]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(mport_o[55]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(mport_o[56]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(mport_o[57]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(mport_o[58]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(mport_o[59]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(mport_o[60]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(mport_o[61]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(mport_o[62]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(mport_o[63]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(mport_o[64]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(mport_o[66]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(mport_o[67]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(pixel_o[0]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(pixel_o[1]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(pixel_o[2]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(pixel_o[3]));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(pixel_o[4]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(pixel_o[5]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(pixel_o[6]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(pixel_o[7]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(vsync_o));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(hsync_o));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(mport_o[34]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(mport_o[35]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(mport_o[36]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(mport_o[37]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(mport_o[38]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(mport_o[39]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(mport_o[40]));
 sky130_fd_sc_hd__conb_1 vga_m_354 (.LO(net354));
 sky130_fd_sc_hd__conb_1 vga_m_355 (.LO(net355));
 sky130_fd_sc_hd__conb_1 vga_m_356 (.LO(net356));
 sky130_fd_sc_hd__conb_1 vga_m_357 (.LO(net357));
 sky130_fd_sc_hd__conb_1 vga_m_358 (.LO(net358));
 sky130_fd_sc_hd__conb_1 vga_m_359 (.LO(net359));
 sky130_fd_sc_hd__conb_1 vga_m_360 (.LO(net360));
 sky130_fd_sc_hd__conb_1 vga_m_361 (.LO(net361));
 sky130_fd_sc_hd__conb_1 vga_m_362 (.LO(net362));
 sky130_fd_sc_hd__conb_1 vga_m_363 (.LO(net363));
 sky130_fd_sc_hd__conb_1 vga_m_364 (.LO(net364));
 sky130_fd_sc_hd__conb_1 vga_m_365 (.LO(net365));
 sky130_fd_sc_hd__conb_1 vga_m_366 (.LO(net366));
 sky130_fd_sc_hd__conb_1 vga_m_367 (.LO(net367));
 sky130_fd_sc_hd__conb_1 vga_m_368 (.LO(net368));
 sky130_fd_sc_hd__conb_1 vga_m_369 (.LO(net369));
 sky130_fd_sc_hd__conb_1 vga_m_370 (.LO(net370));
 sky130_fd_sc_hd__conb_1 vga_m_371 (.LO(net371));
 sky130_fd_sc_hd__conb_1 vga_m_372 (.LO(net372));
 sky130_fd_sc_hd__conb_1 vga_m_373 (.LO(net373));
 sky130_fd_sc_hd__conb_1 vga_m_374 (.LO(net374));
 sky130_fd_sc_hd__conb_1 vga_m_375 (.LO(net375));
 sky130_fd_sc_hd__conb_1 vga_m_376 (.LO(net376));
 sky130_fd_sc_hd__conb_1 vga_m_377 (.LO(net377));
 sky130_fd_sc_hd__conb_1 vga_m_378 (.LO(net378));
 sky130_fd_sc_hd__conb_1 vga_m_379 (.LO(net379));
 sky130_fd_sc_hd__conb_1 vga_m_380 (.LO(net380));
 sky130_fd_sc_hd__conb_1 vga_m_381 (.LO(net381));
 sky130_fd_sc_hd__conb_1 vga_m_382 (.LO(net382));
 sky130_fd_sc_hd__conb_1 vga_m_383 (.LO(net383));
 sky130_fd_sc_hd__conb_1 vga_m_384 (.LO(net384));
 sky130_fd_sc_hd__conb_1 vga_m_385 (.LO(net385));
 sky130_fd_sc_hd__conb_1 vga_m_386 (.LO(net386));
 sky130_fd_sc_hd__conb_1 vga_m_387 (.LO(net387));
 sky130_fd_sc_hd__conb_1 vga_m_388 (.LO(net388));
 sky130_fd_sc_hd__conb_1 vga_m_389 (.LO(net389));
 sky130_fd_sc_hd__buf_6 wire135 (.A(_09495_),
    .X(net135));
 sky130_fd_sc_hd__buf_4 wire136 (.A(_10382_),
    .X(net136));
 assign mport_o[0] = net354;
 assign mport_o[10] = net364;
 assign mport_o[11] = net365;
 assign mport_o[12] = net366;
 assign mport_o[13] = net367;
 assign mport_o[14] = net368;
 assign mport_o[15] = net369;
 assign mport_o[16] = net370;
 assign mport_o[17] = net371;
 assign mport_o[18] = net372;
 assign mport_o[19] = net373;
 assign mport_o[1] = net355;
 assign mport_o[20] = net374;
 assign mport_o[21] = net375;
 assign mport_o[22] = net376;
 assign mport_o[23] = net377;
 assign mport_o[24] = net378;
 assign mport_o[25] = net379;
 assign mport_o[26] = net380;
 assign mport_o[27] = net381;
 assign mport_o[28] = net382;
 assign mport_o[29] = net383;
 assign mport_o[2] = net356;
 assign mport_o[30] = net384;
 assign mport_o[31] = net385;
 assign mport_o[32] = net386;
 assign mport_o[33] = net387;
 assign mport_o[3] = net357;
 assign mport_o[4] = net358;
 assign mport_o[5] = net359;
 assign mport_o[65] = net388;
 assign mport_o[68] = net389;
 assign mport_o[6] = net360;
 assign mport_o[7] = net361;
 assign mport_o[8] = net362;
 assign mport_o[9] = net363;
endmodule

